/opt/tech/tower/digital/tsl18fs190svt_Rev_2019.09/lib/cdl/tsl18fs190svt.cdl