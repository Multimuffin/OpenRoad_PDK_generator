/opt/tech/tower/digital/tsl18fs190svt_Rev_2019.09/lib/lef/tsl18fs190svt.lef