/opt/tech/tower/digital/tsl18fs190svt_Rev_2019.09/tech/lef/3M0L/tsl180l3_0l.lef