
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.6.142
#
# REF LIBS: tsl18fs190svt_wb 
# TECH LIB NAME: ts018_prim
# TECH FILE NAME: techfile.cds
#******

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
    TIME NANOSECONDS 1  ;
    CAPACITANCE PICOFARADS 1  ;
    RESISTANCE OHMS 1  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;
SITE CoreSite
    SYMMETRY Y  ;
    CLASS CORE  ;
    SIZE 0.560 BY 3.920 ;
END CoreSite

MACRO XOR3_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR3_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.775 3.290 2.005 ;
        RECT  2.950 1.260 3.225 2.005 ;
        RECT  1.635 1.260 3.225 1.540 ;
        RECT  1.635 0.435 1.865 1.540 ;
        RECT  0.695 0.435 1.865 0.665 ;
        RECT  0.695 0.435 0.945 1.755 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.670 1.860 4.010 2.465 ;
        RECT  1.760 2.235 4.010 2.465 ;
        RECT  1.390 2.465 2.100 2.760 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.030 1.455 8.870 2.100 ;
        RECT  5.960 1.455 8.870 1.685 ;
        RECT  5.960 1.095 6.190 1.685 ;
        RECT  5.630 1.095 6.190 1.425 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.040 0.470 11.380 3.395 ;
        RECT  9.690 2.695 11.380 3.035 ;
        RECT  11.015 0.700 11.380 3.035 ;
        RECT  9.690 0.700 11.380 1.225 ;
        RECT  9.690 2.695 10.030 3.395 ;
        RECT  9.690 0.470 10.030 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.760 2.575 12.100 4.100 ;
        RECT  8.270 2.890 9.080 4.100 ;
        RECT  6.420 3.110 6.710 4.100 ;
        RECT  1.710 3.110 2.050 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.760 -0.180 12.100 1.345 ;
        RECT  8.970 -0.180 9.310 0.765 ;
        RECT  6.110 -0.180 6.450 0.810 ;
        RECT  3.970 -0.180 4.310 1.150 ;
        RECT  2.095 -0.180 2.380 1.030 ;
        RECT  0.180 -0.180 0.465 1.130 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.175 0.895 1.405 2.235 ;
        RECT  1.175 1.770 2.620 2.005 ;
        RECT  0.480 2.005 1.460 2.235 ;
        RECT  0.480 2.005 0.820 3.295 ;
        RECT  2.470 2.695 2.810 3.450 ;
        RECT  2.470 3.155 4.250 3.450 ;
        RECT  4.775 0.575 5.115 1.885 ;
        RECT  4.775 1.655 5.730 1.885 ;
        RECT  5.445 1.915 6.930 2.200 ;
        RECT  5.445 1.655 5.730 2.975 ;
        RECT  2.760 0.470 3.685 0.810 ;
        RECT  3.455 0.470 3.685 1.610 ;
        RECT  3.455 1.380 4.545 1.610 ;
        RECT  4.315 1.380 4.545 2.925 ;
        RECT  7.160 1.915 7.670 2.200 ;
        RECT  7.160 1.915 7.390 2.660 ;
        RECT  5.960 2.430 7.390 2.660 ;
        RECT  4.315 2.115 5.215 2.925 ;
        RECT  3.190 2.695 5.215 2.925 ;
        RECT  4.920 2.115 5.215 3.510 ;
        RECT  5.960 2.430 6.190 3.510 ;
        RECT  4.920 3.205 6.190 3.510 ;
        RECT  6.830 0.470 8.610 0.765 ;
        RECT  6.830 0.470 7.170 1.225 ;
        RECT  7.550 0.995 9.460 1.225 ;
        RECT  9.230 1.620 10.675 1.960 ;
        RECT  9.230 0.995 9.460 2.660 ;
        RECT  7.620 2.430 9.460 2.660 ;
        RECT  7.620 2.430 7.850 3.450 ;
        RECT  7.090 3.110 7.850 3.450 ;
    END
END XOR3_X8_18_SVT_WB

MACRO XOR3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.875 1.235 3.160 1.960 ;
        RECT  1.530 1.235 3.160 1.465 ;
        RECT  1.530 0.410 1.760 1.465 ;
        RECT  0.130 0.410 1.760 0.640 ;
        RECT  0.130 1.270 0.840 1.730 ;
        RECT  0.130 0.410 0.465 1.730 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.575 1.915 3.915 2.420 ;
        RECT  1.760 2.190 3.915 2.420 ;
        RECT  1.295 2.420 2.100 2.760 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.740 1.455 8.550 1.960 ;
        RECT  5.765 1.455 8.550 1.685 ;
        RECT  5.460 1.160 6.140 1.540 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.400 2.470 10.525 2.700 ;
        RECT  10.200 1.440 10.525 2.700 ;
        RECT  9.400 1.440 10.525 1.670 ;
        RECT  9.400 2.470 9.940 3.395 ;
        RECT  9.400 0.685 9.740 1.670 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  10.170 3.110 10.460 4.100 ;
        RECT  7.980 3.110 8.790 4.100 ;
        RECT  6.165 3.100 6.450 4.100 ;
        RECT  1.655 3.110 1.995 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  10.120 -0.180 10.460 1.210 ;
        RECT  8.680 -0.180 9.020 0.765 ;
        RECT  5.780 -0.180 6.120 0.915 ;
        RECT  3.850 -0.180 4.190 1.225 ;
        RECT  1.990 -0.180 2.275 1.005 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.070 1.695 2.495 1.960 ;
        RECT  1.070 0.870 1.300 2.190 ;
        RECT  0.385 1.960 1.300 2.190 ;
        RECT  0.385 1.960 0.725 3.295 ;
        RECT  2.375 2.650 2.715 3.450 ;
        RECT  2.375 3.110 4.155 3.450 ;
        RECT  4.605 0.575 5.230 1.540 ;
        RECT  5.000 0.575 5.230 2.720 ;
        RECT  5.000 1.915 6.670 2.190 ;
        RECT  5.000 1.915 5.475 2.720 ;
        RECT  2.655 0.660 3.620 1.000 ;
        RECT  3.390 0.660 3.620 1.685 ;
        RECT  3.390 1.455 4.375 1.685 ;
        RECT  4.145 1.455 4.375 2.880 ;
        RECT  6.900 1.915 7.410 2.200 ;
        RECT  6.900 1.915 7.130 2.650 ;
        RECT  5.705 2.420 7.130 2.650 ;
        RECT  4.145 1.915 4.670 2.880 ;
        RECT  3.095 2.650 4.670 2.880 ;
        RECT  4.385 1.915 4.670 3.290 ;
        RECT  5.705 2.420 5.935 3.290 ;
        RECT  4.385 2.950 5.935 3.290 ;
        RECT  6.540 0.470 8.320 0.765 ;
        RECT  6.540 0.470 6.880 1.225 ;
        RECT  7.260 0.995 9.170 1.225 ;
        RECT  8.940 1.900 9.970 2.200 ;
        RECT  7.360 2.540 9.170 2.880 ;
        RECT  8.940 0.995 9.170 2.880 ;
        RECT  6.830 2.880 7.590 3.220 ;
    END
END XOR3_X4_18_SVT_WB

MACRO XOR3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.380 3.140 2.725 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.760 3.950 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.920 1.915 8.260 2.400 ;
        RECT  5.980 2.170 8.260 2.400 ;
        RECT  5.690 2.380 6.310 2.695 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.700 2.630 8.820 2.870 ;
        RECT  8.520 1.455 8.820 2.870 ;
        RECT  7.770 1.455 8.820 1.685 ;
        RECT  7.770 0.470 8.000 1.685 ;
        RECT  6.980 0.470 8.000 0.810 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  6.220 3.045 6.560 4.100 ;
        RECT  1.850 3.015 2.190 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.420 -0.180 8.760 1.225 ;
        RECT  4.130 -0.180 4.470 0.695 ;
        RECT  1.850 -0.180 2.190 0.925 ;
        RECT  0.330 -0.180 0.670 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.090 0.640 1.430 1.500 ;
        RECT  0.230 1.160 2.380 1.500 ;
        RECT  0.230 1.160 0.595 3.295 ;
        RECT  0.230 2.955 0.945 3.295 ;
        RECT  2.610 3.055 2.950 3.395 ;
        RECT  4.090 2.790 4.430 3.395 ;
        RECT  2.610 3.150 4.430 3.395 ;
        RECT  5.265 0.925 5.800 1.940 ;
        RECT  5.265 1.640 6.840 1.940 ;
        RECT  5.265 0.925 5.495 2.245 ;
        RECT  4.790 2.015 5.495 2.245 ;
        RECT  4.790 2.015 5.130 3.395 ;
        RECT  4.805 0.410 6.370 0.695 ;
        RECT  2.610 0.695 3.710 1.175 ;
        RECT  2.610 0.945 5.035 1.175 ;
        RECT  6.030 0.410 6.370 1.410 ;
        RECT  6.030 1.180 7.540 1.410 ;
        RECT  4.805 0.410 5.035 1.785 ;
        RECT  4.280 0.945 5.035 1.785 ;
        RECT  7.200 1.180 7.540 1.940 ;
        RECT  4.280 0.945 4.560 2.560 ;
        RECT  3.370 2.330 4.560 2.560 ;
        RECT  3.370 2.330 3.710 2.920 ;
        RECT  6.980 2.630 7.320 3.385 ;
        RECT  6.980 3.100 8.760 3.385 ;
    END
END XOR3_X2_18_SVT_WB

MACRO XOR3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.375 2.030 2.885 2.325 ;
        RECT  0.650 2.380 2.605 2.815 ;
        RECT  2.375 2.030 2.605 2.815 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.280 1.570 3.620 2.275 ;
        RECT  0.970 1.570 3.620 1.800 ;
        RECT  0.970 1.570 1.620 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.730 1.720 7.720 2.150 ;
        RECT  5.490 2.480 6.960 2.770 ;
        RECT  6.730 1.720 6.960 2.770 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.687  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.190 2.380 8.285 2.610 ;
        RECT  7.950 0.585 8.285 2.610 ;
        RECT  6.690 0.585 8.285 0.875 ;
        RECT  7.190 2.380 7.500 2.970 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  5.680 3.000 6.020 4.100 ;
        RECT  1.560 3.045 1.900 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.880 -0.180 8.220 0.355 ;
        RECT  3.800 -0.180 4.140 0.820 ;
        RECT  1.560 -0.180 1.900 0.820 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.800 0.535 1.140 1.340 ;
        RECT  0.190 1.055 2.075 1.340 ;
        RECT  0.190 1.055 0.420 3.385 ;
        RECT  0.190 3.045 0.710 3.385 ;
        RECT  4.835 1.005 5.535 2.250 ;
        RECT  4.835 2.010 6.500 2.250 ;
        RECT  4.530 2.095 5.010 3.290 ;
        RECT  4.370 0.545 6.425 0.775 ;
        RECT  2.320 0.535 2.660 1.280 ;
        RECT  6.160 0.545 6.425 1.445 ;
        RECT  2.320 1.050 4.605 1.280 ;
        RECT  6.160 1.105 7.250 1.445 ;
        RECT  4.370 0.545 4.605 1.865 ;
        RECT  3.850 1.050 4.605 1.865 ;
        RECT  3.850 1.050 4.080 2.845 ;
        RECT  3.040 2.505 4.080 2.845 ;
        RECT  6.400 3.105 6.740 3.445 ;
        RECT  7.880 2.840 8.220 3.445 ;
        RECT  6.400 3.215 8.220 3.445 ;
    END
END XOR3_X1_18_SVT_WB

MACRO XOR3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.490 2.085 3.000 2.380 ;
        RECT  0.715 2.380 2.720 2.720 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.380 1.625 3.720 1.920 ;
        RECT  1.260 1.625 3.720 1.855 ;
        RECT  1.260 1.625 1.720 2.150 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.390 1.625 7.730 2.190 ;
        RECT  5.500 1.625 7.730 1.855 ;
        RECT  5.500 1.625 5.860 2.150 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.150 2.570 8.260 2.910 ;
        RECT  7.960 1.105 8.260 2.910 ;
        RECT  7.235 1.105 8.260 1.395 ;
        RECT  7.235 0.535 7.580 1.395 ;
        RECT  6.430 0.535 7.580 0.825 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  5.615 3.350 5.955 4.100 ;
        RECT  1.620 2.990 1.960 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.870 -0.180 8.210 0.875 ;
        RECT  3.860 -0.180 4.200 0.875 ;
        RECT  1.660 -0.180 2.000 0.825 ;
        RECT  0.180 -0.180 0.520 0.825 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.535 1.240 1.395 ;
        RECT  0.180 1.055 2.190 1.395 ;
        RECT  0.180 1.055 0.485 3.330 ;
        RECT  4.980 0.535 5.320 1.395 ;
        RECT  4.410 1.055 5.320 1.395 ;
        RECT  4.410 1.105 6.295 1.395 ;
        RECT  4.410 1.055 4.640 2.910 ;
        RECT  4.410 2.570 4.810 2.910 ;
        RECT  2.420 0.535 2.760 1.395 ;
        RECT  2.420 1.105 4.180 1.395 ;
        RECT  4.870 1.780 5.270 2.335 ;
        RECT  5.040 1.780 5.270 3.510 ;
        RECT  6.500 2.085 7.010 2.380 ;
        RECT  5.040 2.380 6.730 2.720 ;
        RECT  3.140 2.570 4.180 2.910 ;
        RECT  3.950 1.105 4.180 3.510 ;
        RECT  5.040 2.380 5.340 3.510 ;
        RECT  3.950 3.255 5.340 3.510 ;
    END
END XOR3_X0_18_SVT_WB

MACRO XOR2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.680 1.915 3.190 2.200 ;
        RECT  1.490 2.380 2.910 2.660 ;
        RECT  2.680 1.915 2.910 2.660 ;
        RECT  0.515 3.160 1.720 3.390 ;
        RECT  1.490 2.380 1.720 3.390 ;
        RECT  0.515 2.070 0.800 3.390 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.540 1.455 4.350 2.150 ;
        RECT  1.545 1.455 4.350 1.685 ;
        RECT  1.545 1.095 1.775 1.685 ;
        RECT  1.260 1.095 1.775 1.380 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.505 2.250 7.000 3.135 ;
        RECT  6.770 0.650 7.000 3.135 ;
        RECT  5.065 1.050 7.000 1.390 ;
        RECT  6.300 0.650 7.000 1.390 ;
        RECT  5.065 2.250 7.000 2.480 ;
        RECT  5.065 2.250 5.405 3.135 ;
        RECT  5.065 0.660 5.405 1.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  7.230 2.575 7.570 4.100 ;
        RECT  5.785 2.710 6.125 4.100 ;
        RECT  3.780 3.070 4.590 4.100 ;
        RECT  1.925 3.515 2.210 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  7.230 -0.180 7.570 1.290 ;
        RECT  5.785 -0.180 6.070 0.810 ;
        RECT  1.580 -0.180 1.920 0.865 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.350 0.575 0.690 1.840 ;
        RECT  0.350 1.610 1.315 1.840 ;
        RECT  1.030 1.610 1.315 2.150 ;
        RECT  1.030 1.915 2.450 2.150 ;
        RECT  1.030 1.610 1.260 2.930 ;
        RECT  2.340 0.470 4.120 0.765 ;
        RECT  3.060 0.995 4.810 1.225 ;
        RECT  4.580 1.620 6.540 1.960 ;
        RECT  4.580 0.995 4.810 2.785 ;
        RECT  3.140 2.445 4.810 2.785 ;
        RECT  3.140 2.445 3.370 3.185 ;
        RECT  2.630 2.890 3.370 3.185 ;
    END
END XOR2_X8_18_SVT_WB

MACRO XOR2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.690 2.380 3.385 2.660 ;
        RECT  3.045 1.915 3.385 2.660 ;
        RECT  0.740 3.160 1.920 3.500 ;
        RECT  1.690 2.380 1.920 3.500 ;
        RECT  0.740 2.070 1.000 3.500 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.765 1.455 4.575 2.100 ;
        RECT  1.765 1.455 4.575 1.685 ;
        RECT  1.765 1.095 1.995 1.685 ;
        RECT  1.485 1.095 1.995 1.380 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.740 1.065 6.020 2.705 ;
        RECT  5.465 2.430 5.805 3.185 ;
        RECT  5.465 0.675 5.805 1.405 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  6.250 2.660 6.535 4.100 ;
        RECT  4.235 3.045 5.045 4.100 ;
        RECT  2.150 2.890 2.435 4.100 ;
        RECT  0.195 2.590 0.510 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.250 -0.180 6.535 1.255 ;
        RECT  4.705 -0.180 5.045 0.490 ;
        RECT  1.805 -0.180 2.145 0.865 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.575 0.575 0.915 1.840 ;
        RECT  0.575 1.610 1.515 1.840 ;
        RECT  1.230 1.610 1.515 2.150 ;
        RECT  1.230 1.915 2.685 2.150 ;
        RECT  1.230 1.610 1.460 2.930 ;
        RECT  2.565 0.470 4.345 0.765 ;
        RECT  3.285 0.995 5.200 1.225 ;
        RECT  4.860 1.860 5.510 2.200 ;
        RECT  4.860 0.995 5.200 2.670 ;
        RECT  3.615 2.330 5.200 2.670 ;
        RECT  3.615 2.330 3.845 3.405 ;
        RECT  2.855 3.065 3.845 3.405 ;
    END
END XOR2_X4_18_SVT_WB

MACRO XOR2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.895 1.915 3.405 2.180 ;
        RECT  1.680 2.375 3.125 2.655 ;
        RECT  2.895 1.915 3.125 2.655 ;
        RECT  0.700 3.270 1.910 3.500 ;
        RECT  1.680 2.375 1.910 3.500 ;
        RECT  0.700 2.180 0.990 3.500 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.755 1.455 4.565 2.100 ;
        RECT  1.755 1.455 4.565 1.685 ;
        RECT  1.475 1.160 1.985 1.455 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.888  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.415 2.390 6.550 2.620 ;
        RECT  6.215 1.105 6.550 2.620 ;
        RECT  5.415 1.105 6.550 1.335 ;
        RECT  5.415 2.390 6.020 3.270 ;
        RECT  5.415 0.810 5.755 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  6.250 2.850 6.535 4.100 ;
        RECT  4.035 3.430 4.845 4.100 ;
        RECT  2.140 2.920 2.425 4.100 ;
        RECT  0.185 2.740 0.470 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.175 -0.180 6.515 0.875 ;
        RECT  4.695 -0.180 5.035 0.765 ;
        RECT  1.795 -0.180 2.135 0.915 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.565 0.575 0.905 1.915 ;
        RECT  0.565 1.685 1.505 1.915 ;
        RECT  1.220 1.915 2.665 2.145 ;
        RECT  1.220 1.685 1.450 3.040 ;
        RECT  2.555 0.470 4.335 0.765 ;
        RECT  2.555 0.470 2.895 1.225 ;
        RECT  3.275 0.995 5.185 1.225 ;
        RECT  4.900 1.840 5.985 2.160 ;
        RECT  4.900 0.995 5.185 3.195 ;
        RECT  2.845 2.885 5.185 3.195 ;
    END
END XOR2_X3_18_SVT_WB

MACRO XOR2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.630 3.430 1.970 ;
        RECT  2.920 1.280 3.150 1.970 ;
        RECT  1.670 1.280 3.150 1.510 ;
        RECT  1.670 0.410 1.900 1.510 ;
        RECT  0.700 0.410 1.900 0.640 ;
        RECT  0.700 0.410 0.980 1.730 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.790 1.860 4.130 2.430 ;
        RECT  1.790 2.200 4.130 2.430 ;
        RECT  1.510 2.430 2.100 2.770 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.310 2.660 4.900 2.890 ;
        RECT  4.560 1.035 4.900 2.890 ;
        RECT  3.440 1.035 4.900 1.375 ;
        RECT  3.440 0.500 3.780 1.375 ;
        RECT  2.850 0.500 3.780 0.840 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  1.870 3.000 2.210 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.030 -0.180 4.370 0.805 ;
        RECT  2.130 -0.180 2.470 1.050 ;
        RECT  0.185 -0.180 0.470 1.105 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.210 0.870 1.440 2.200 ;
        RECT  1.210 1.740 2.690 1.970 ;
        RECT  0.600 1.970 1.550 2.200 ;
        RECT  0.600 1.970 0.940 3.385 ;
        RECT  2.590 3.120 4.370 3.450 ;
    END
END XOR2_X2_18_SVT_WB

MACRO XOR2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.670 2.375 2.950 2.715 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.770 3.740 2.125 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.687  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.180 2.385 4.270 2.615 ;
        RECT  3.970 1.200 4.270 2.615 ;
        RECT  3.180 1.200 4.270 1.540 ;
        RECT  3.180 2.385 3.520 2.975 ;
        RECT  3.180 0.590 3.520 1.540 ;
        RECT  2.420 0.590 3.520 0.930 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  1.660 2.955 2.000 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.940 -0.180 4.280 0.930 ;
        RECT  1.660 -0.180 2.000 0.875 ;
        RECT  0.180 -0.180 0.520 0.880 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.590 1.240 1.450 ;
        RECT  0.190 1.110 2.200 1.450 ;
        RECT  0.190 1.110 0.420 3.295 ;
        RECT  0.190 2.955 0.810 3.295 ;
        RECT  2.420 3.110 2.760 3.450 ;
        RECT  3.900 2.845 4.240 3.450 ;
        RECT  2.420 3.205 4.240 3.450 ;
    END
END XOR2_X1_18_SVT_WB

MACRO XOR2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.440 2.090 2.950 2.375 ;
        RECT  0.715 2.380 2.670 2.720 ;
        RECT  2.440 2.090 2.670 2.720 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.400 1.565 3.740 1.905 ;
        RECT  1.210 1.630 3.740 1.860 ;
        RECT  1.210 1.630 1.720 2.100 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.462  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.160 2.595 4.340 3.020 ;
        RECT  4.000 1.055 4.340 3.020 ;
        RECT  2.420 1.055 4.340 1.335 ;
        RECT  2.420 0.540 2.760 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  1.700 2.975 2.040 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.880 -0.180 4.220 0.825 ;
        RECT  1.660 -0.180 2.000 0.830 ;
        RECT  0.180 -0.180 0.520 0.830 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.540 1.240 1.400 ;
        RECT  0.180 1.060 2.190 1.400 ;
        RECT  0.180 1.060 0.485 3.315 ;
    END
END XOR2_X0_18_SVT_WB

MACRO XOR2NG_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2NG_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.285 1.595 3.780 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.910 0.760 2.200 ;
        RECT  0.140 1.910 0.480 2.765 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.620 2.130 2.585 2.360 ;
        RECT  2.355 0.990 2.585 2.360 ;
        RECT  2.050 0.990 2.585 1.330 ;
        RECT  1.620 2.130 2.100 2.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.050 3.460 3.440 4.100 ;
        RECT  0.220 3.460 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.400 -0.180 3.740 0.460 ;
        RECT  0.900 -0.180 1.240 1.220 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.040 0.520 1.680 ;
        RECT  0.180 1.450 1.330 1.680 ;
        RECT  0.990 1.560 2.125 1.900 ;
        RECT  0.990 1.450 1.240 2.855 ;
        RECT  0.900 2.515 1.240 2.855 ;
        RECT  2.815 1.040 3.055 2.930 ;
        RECT  2.340 2.590 3.055 2.930 ;
        RECT  2.340 2.590 2.680 3.395 ;
        RECT  1.380 3.055 2.680 3.395 ;
    END
END XOR2NG_X1_18_SVT_WB

MACRO XOR2NG_X1P5_18_SVT_WB
    CLASS CORE ;
    FOREIGN XOR2NG_X1P5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.335  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.325 1.770 3.805 2.195 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.915 0.800 2.200 ;
        RECT  0.140 1.915 0.480 2.710 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.643  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.660 2.220 2.625 2.450 ;
        RECT  2.395 0.995 2.625 2.450 ;
        RECT  2.100 0.995 2.625 1.335 ;
        RECT  1.660 2.220 2.100 2.745 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.140 3.460 3.480 4.100 ;
        RECT  0.180 3.460 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.400 -0.180 3.740 0.405 ;
        RECT  0.940 -0.180 1.280 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.045 0.560 1.685 ;
        RECT  0.220 1.455 1.370 1.685 ;
        RECT  1.030 1.565 2.165 1.905 ;
        RECT  1.030 1.455 1.280 2.965 ;
        RECT  0.940 2.625 1.280 2.965 ;
        RECT  2.855 1.045 3.095 3.020 ;
        RECT  2.380 2.680 3.095 3.020 ;
        RECT  2.380 2.680 2.720 3.485 ;
        RECT  1.425 3.145 2.720 3.485 ;
    END
END XOR2NG_X1P5_18_SVT_WB

MACRO XNOR3_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR3_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.050 1.235 3.390 1.960 ;
        RECT  1.590 1.235 3.390 1.465 ;
        RECT  1.590 0.640 1.895 1.465 ;
        RECT  0.140 0.640 1.895 0.870 ;
        RECT  0.140 1.620 0.845 1.960 ;
        RECT  0.140 0.640 0.480 1.960 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.535 2.200 4.075 2.430 ;
        RECT  3.770 1.860 4.075 2.430 ;
        RECT  1.535 2.200 2.100 2.770 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.665 2.165 8.830 2.395 ;
        RECT  8.020 1.770 8.830 2.395 ;
        RECT  5.665 2.165 6.080 2.505 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.680 1.040 11.620 1.280 ;
        RECT  11.120 0.525 11.620 1.280 ;
        RECT  11.120 0.525 11.460 3.395 ;
        RECT  9.680 2.250 11.460 2.480 ;
        RECT  9.680 2.250 10.020 3.170 ;
        RECT  9.680 0.525 10.020 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  10.400 2.710 10.740 4.100 ;
        RECT  8.960 3.150 9.300 4.100 ;
        RECT  6.100 3.105 6.440 4.100 ;
        RECT  1.850 3.105 2.190 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  10.400 -0.180 10.740 0.810 ;
        RECT  8.260 -0.180 9.070 0.810 ;
        RECT  6.380 -0.180 6.720 0.810 ;
        RECT  4.080 -0.180 4.420 1.170 ;
        RECT  2.125 -0.180 2.400 0.930 ;
        RECT  0.180 -0.180 2.400 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.075 1.100 1.360 1.970 ;
        RECT  1.075 1.695 2.690 1.970 ;
        RECT  1.075 1.100 1.305 2.430 ;
        RECT  0.580 2.200 1.305 2.430 ;
        RECT  0.580 2.200 0.920 3.295 ;
        RECT  2.570 2.690 2.910 3.445 ;
        RECT  2.570 3.150 4.350 3.445 ;
        RECT  5.195 0.995 5.490 1.935 ;
        RECT  5.195 1.620 6.920 1.935 ;
        RECT  5.195 0.995 5.435 3.295 ;
        RECT  4.765 2.690 5.435 3.295 ;
        RECT  4.680 0.425 6.060 0.765 ;
        RECT  2.830 0.590 3.850 0.930 ;
        RECT  5.720 0.425 6.060 1.390 ;
        RECT  5.720 1.050 7.380 1.390 ;
        RECT  3.620 0.590 3.850 1.630 ;
        RECT  7.150 1.050 7.380 1.935 ;
        RECT  3.620 1.400 4.965 1.630 ;
        RECT  7.150 1.620 7.660 1.935 ;
        RECT  4.680 0.425 4.965 2.430 ;
        RECT  4.305 1.400 4.965 2.430 ;
        RECT  4.305 1.400 4.535 2.920 ;
        RECT  3.290 2.660 4.535 2.920 ;
        RECT  6.820 2.690 7.160 3.445 ;
        RECT  6.820 3.150 8.600 3.445 ;
        RECT  7.100 0.470 7.840 0.810 ;
        RECT  7.610 0.470 7.840 1.380 ;
        RECT  7.610 1.040 9.450 1.380 ;
        RECT  9.220 1.620 10.665 1.960 ;
        RECT  9.220 1.040 9.450 2.920 ;
        RECT  7.540 2.635 9.450 2.920 ;
    END
END XNOR3_X8_18_SVT_WB

MACRO XNOR3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.020 1.770 3.530 2.000 ;
        RECT  3.020 1.160 3.250 2.000 ;
        RECT  1.845 1.160 3.250 1.390 ;
        RECT  1.845 0.640 2.075 1.390 ;
        RECT  0.140 0.640 2.075 0.870 ;
        RECT  0.140 1.670 0.960 1.955 ;
        RECT  0.140 0.640 0.495 1.955 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.650 2.230 4.185 2.460 ;
        RECT  3.880 1.860 4.185 2.460 ;
        RECT  1.650 2.230 2.100 2.755 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.130 1.860 8.940 2.420 ;
        RECT  6.240 2.190 8.940 2.420 ;
        RECT  5.785 2.415 6.580 2.755 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.090 0.590 10.320 2.555 ;
        RECT  9.790 2.325 10.130 3.175 ;
        RECT  9.660 0.590 10.320 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  10.510 2.695 10.850 4.100 ;
        RECT  9.070 3.165 9.410 4.100 ;
        RECT  6.210 3.110 6.550 4.100 ;
        RECT  1.960 3.110 2.300 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  10.550 -0.180 10.890 1.165 ;
        RECT  8.370 -0.180 9.180 0.810 ;
        RECT  6.490 -0.180 6.830 0.820 ;
        RECT  4.160 -0.180 4.500 1.125 ;
        RECT  2.305 -0.180 2.535 0.930 ;
        RECT  0.225 -0.180 2.535 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.860 1.100 1.615 1.440 ;
        RECT  1.190 1.100 1.615 1.960 ;
        RECT  1.190 1.620 2.790 1.960 ;
        RECT  1.190 1.100 1.420 2.475 ;
        RECT  0.220 2.185 1.420 2.475 ;
        RECT  0.220 2.185 1.030 3.450 ;
        RECT  2.680 2.690 3.020 3.445 ;
        RECT  2.680 3.150 4.460 3.445 ;
        RECT  5.315 0.995 5.610 1.960 ;
        RECT  5.315 1.730 7.050 1.960 ;
        RECT  5.315 0.995 5.555 2.835 ;
        RECT  4.875 2.590 5.555 2.835 ;
        RECT  4.875 2.590 5.160 3.295 ;
        RECT  4.800 0.425 6.180 0.765 ;
        RECT  2.970 0.540 3.905 0.880 ;
        RECT  5.840 0.425 6.180 1.500 ;
        RECT  3.675 0.540 3.905 1.585 ;
        RECT  5.840 1.270 7.510 1.500 ;
        RECT  3.675 1.355 5.085 1.585 ;
        RECT  7.280 1.270 7.510 1.960 ;
        RECT  7.280 1.620 7.790 1.960 ;
        RECT  4.800 0.425 5.085 1.980 ;
        RECT  4.415 1.355 5.085 1.980 ;
        RECT  4.415 1.355 4.645 2.920 ;
        RECT  3.400 2.690 4.645 2.920 ;
        RECT  6.930 2.690 7.270 3.445 ;
        RECT  6.930 3.165 8.710 3.445 ;
        RECT  7.210 0.700 7.970 1.040 ;
        RECT  7.740 1.040 9.430 1.380 ;
        RECT  9.200 1.040 9.430 2.935 ;
        RECT  9.200 1.620 9.860 1.960 ;
        RECT  9.200 1.620 9.540 2.935 ;
        RECT  7.650 2.650 9.540 2.935 ;
    END
END XNOR3_X4_18_SVT_WB

MACRO XNOR3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.730 2.380 2.990 2.775 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.820 3.780 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.090 1.455 8.385 1.960 ;
        RECT  5.975 1.455 8.385 1.685 ;
        RECT  5.975 1.160 6.580 1.685 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.910 2.330 8.845 2.710 ;
        RECT  8.615 0.985 8.845 2.710 ;
        RECT  7.720 0.985 8.845 1.225 ;
        RECT  7.180 3.110 8.140 3.450 ;
        RECT  7.910 2.330 8.140 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.370 2.990 8.710 4.100 ;
        RECT  4.010 3.570 4.820 4.100 ;
        RECT  1.700 3.015 2.040 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  6.240 -0.180 6.580 0.915 ;
        RECT  3.940 -0.180 4.280 0.820 ;
        RECT  1.700 -0.180 2.040 0.935 ;
        RECT  0.180 -0.180 0.520 0.940 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.650 1.280 1.510 ;
        RECT  0.270 1.170 2.240 1.510 ;
        RECT  0.270 1.170 0.500 3.295 ;
        RECT  0.270 3.005 0.850 3.295 ;
        RECT  2.460 3.055 2.800 3.340 ;
        RECT  3.940 2.790 4.280 3.340 ;
        RECT  2.460 3.110 4.280 3.340 ;
        RECT  5.065 0.535 5.350 1.045 ;
        RECT  5.065 0.815 5.745 1.045 ;
        RECT  5.515 0.815 5.745 2.720 ;
        RECT  5.515 1.915 7.020 2.200 ;
        RECT  5.515 1.915 6.020 2.720 ;
        RECT  2.460 0.650 3.080 0.990 ;
        RECT  2.740 0.650 3.080 1.590 ;
        RECT  2.740 1.250 4.940 1.590 ;
        RECT  7.250 1.915 7.760 2.150 ;
        RECT  4.940 1.360 5.285 2.560 ;
        RECT  3.220 2.330 5.285 2.560 ;
        RECT  7.250 1.915 7.480 2.770 ;
        RECT  6.250 2.430 7.480 2.770 ;
        RECT  3.220 2.330 3.560 2.880 ;
        RECT  5.000 1.360 5.285 3.290 ;
        RECT  6.250 2.430 6.590 3.290 ;
        RECT  5.000 2.950 6.590 3.290 ;
        RECT  7.000 0.470 8.780 0.755 ;
        RECT  7.000 0.470 7.340 1.225 ;
    END
END XNOR3_X2_18_SVT_WB

MACRO XNOR3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.505 2.030 3.015 2.325 ;
        RECT  0.730 2.380 2.735 2.815 ;
        RECT  2.505 2.030 2.735 2.815 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.350 1.570 3.780 2.275 ;
        RECT  1.410 1.570 3.780 1.800 ;
        RECT  1.410 1.570 1.830 2.065 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.660 1.945 8.260 2.175 ;
        RECT  7.920 1.770 8.260 2.175 ;
        RECT  5.660 1.945 6.000 2.410 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.240 2.440 8.810 2.780 ;
        RECT  8.490 1.265 8.810 2.780 ;
        RECT  7.680 1.265 8.810 1.495 ;
        RECT  7.680 0.910 8.020 1.495 ;
        RECT  6.860 2.865 7.470 3.270 ;
        RECT  7.240 2.440 7.470 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.440 3.055 8.780 4.100 ;
        RECT  6.200 3.400 6.540 4.100 ;
        RECT  4.650 3.100 4.990 4.100 ;
        RECT  1.640 3.045 1.980 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  6.200 -0.180 6.540 0.820 ;
        RECT  1.680 -0.180 2.020 0.820 ;
        RECT  0.200 -0.180 0.540 0.825 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.920 0.535 1.260 1.340 ;
        RECT  0.200 1.055 2.220 1.340 ;
        RECT  0.200 1.055 0.500 3.385 ;
        RECT  4.540 0.870 5.350 1.145 ;
        RECT  6.230 2.405 6.740 2.635 ;
        RECT  4.540 0.870 4.770 2.870 ;
        RECT  6.230 2.405 6.460 2.870 ;
        RECT  4.540 2.640 6.460 2.870 ;
        RECT  5.440 2.640 5.780 3.265 ;
        RECT  2.480 0.535 2.780 0.895 ;
        RECT  4.010 0.410 5.920 0.640 ;
        RECT  2.480 0.605 4.240 0.895 ;
        RECT  5.580 0.410 5.920 1.715 ;
        RECT  5.170 1.375 7.450 1.715 ;
        RECT  4.010 0.410 4.240 2.845 ;
        RECT  3.165 2.505 4.240 2.845 ;
        RECT  6.960 0.450 8.740 0.680 ;
        RECT  8.400 0.450 8.740 1.035 ;
        RECT  6.960 0.450 7.300 1.145 ;
    END
END XNOR3_X1_18_SVT_WB

MACRO XNOR3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.510 2.040 3.020 2.325 ;
        RECT  0.735 2.380 2.740 2.720 ;
        RECT  2.510 2.040 2.740 2.720 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.400 1.515 3.740 1.855 ;
        RECT  1.260 1.580 3.740 1.810 ;
        RECT  1.260 1.580 1.740 2.150 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.765 2.120 8.265 2.350 ;
        RECT  7.945 1.765 8.265 2.350 ;
        RECT  5.765 1.895 6.140 2.350 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.820 2.580 8.820 2.815 ;
        RECT  8.520 1.075 8.820 2.815 ;
        RECT  7.550 1.075 8.820 1.415 ;
        RECT  6.820 2.580 7.160 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.260 3.045 8.600 4.100 ;
        RECT  6.060 3.095 6.400 4.100 ;
        RECT  4.580 3.095 4.920 4.100 ;
        RECT  1.640 3.045 1.980 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  6.020 -0.180 6.360 1.155 ;
        RECT  1.680 -0.180 2.020 0.825 ;
        RECT  0.200 -0.180 0.540 0.825 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.920 0.535 1.260 1.350 ;
        RECT  0.200 1.055 2.210 1.350 ;
        RECT  0.200 1.055 0.505 3.385 ;
        RECT  4.580 0.870 4.885 2.865 ;
        RECT  4.580 2.580 6.590 2.865 ;
        RECT  5.300 2.580 5.640 3.385 ;
        RECT  4.000 0.410 5.395 0.640 ;
        RECT  2.440 0.535 2.780 1.285 ;
        RECT  2.440 1.055 4.285 1.285 ;
        RECT  5.115 1.385 7.120 1.665 ;
        RECT  6.890 1.595 7.400 1.890 ;
        RECT  5.115 0.410 5.395 2.180 ;
        RECT  4.000 0.410 4.285 2.845 ;
        RECT  3.170 2.505 4.285 2.845 ;
    END
END XNOR3_X0_18_SVT_WB

MACRO XNOR2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.165 3.220 1.905 ;
        RECT  1.530 1.165 3.220 1.420 ;
        RECT  1.530 0.580 1.760 1.420 ;
        RECT  0.445 0.580 1.760 0.810 ;
        RECT  0.445 1.535 0.840 1.790 ;
        RECT  0.445 0.580 0.675 1.790 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.530 2.135 4.380 2.365 ;
        RECT  3.570 1.760 4.380 2.365 ;
        RECT  1.170 2.480 1.760 2.775 ;
        RECT  1.530 2.135 1.760 2.775 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.670 0.525 7.140 1.590 ;
        RECT  6.670 0.525 7.010 3.395 ;
        RECT  5.230 2.640 7.010 2.880 ;
        RECT  6.660 1.040 7.010 2.880 ;
        RECT  5.230 1.040 7.140 1.350 ;
        RECT  5.230 2.640 5.570 3.395 ;
        RECT  5.230 0.595 5.570 1.350 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.950 3.110 6.290 4.100 ;
        RECT  4.510 3.110 4.850 4.100 ;
        RECT  1.650 3.110 1.990 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.950 -0.180 6.290 0.810 ;
        RECT  3.895 -0.180 4.705 0.410 ;
        RECT  1.990 -0.180 2.280 0.855 ;
        RECT  0.185 -0.180 2.280 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.905 1.040 1.300 1.305 ;
        RECT  1.070 1.650 2.520 1.905 ;
        RECT  1.070 1.040 1.300 2.250 ;
        RECT  0.260 2.020 1.300 2.250 ;
        RECT  0.260 2.020 0.600 3.295 ;
        RECT  2.370 3.110 4.150 3.450 ;
        RECT  2.660 0.650 5.000 0.935 ;
        RECT  4.695 1.620 5.985 1.960 ;
        RECT  4.695 0.650 5.000 2.880 ;
        RECT  3.090 2.595 5.000 2.880 ;
    END
END XNOR2_X8_18_SVT_WB

MACRO XNOR2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.100 1.200 3.440 1.960 ;
        RECT  1.735 1.200 3.440 1.540 ;
        RECT  1.735 0.580 1.965 1.540 ;
        RECT  0.700 0.580 1.965 0.815 ;
        RECT  0.700 1.535 1.045 1.795 ;
        RECT  0.700 0.580 0.930 1.795 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.735 2.230 4.610 2.460 ;
        RECT  3.800 1.820 4.610 2.460 ;
        RECT  1.400 2.485 1.965 2.775 ;
        RECT  1.735 2.230 1.965 2.775 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.770 0.470 6.020 2.480 ;
        RECT  5.475 2.245 5.785 3.230 ;
        RECT  5.450 0.470 6.020 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  6.195 2.695 6.535 4.100 ;
        RECT  4.755 3.165 5.095 4.100 ;
        RECT  1.880 3.110 2.220 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.250 -0.180 6.535 1.305 ;
        RECT  4.080 -0.180 4.890 0.410 ;
        RECT  2.195 -0.180 2.445 0.875 ;
        RECT  0.185 -0.180 2.445 0.350 ;
        RECT  0.185 -0.180 0.470 0.905 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.160 1.045 1.505 1.320 ;
        RECT  1.275 1.770 2.720 2.000 ;
        RECT  1.275 1.045 1.505 2.255 ;
        RECT  0.490 2.025 1.505 2.255 ;
        RECT  0.490 2.025 0.830 3.295 ;
        RECT  2.600 2.690 2.940 3.445 ;
        RECT  2.600 3.165 4.380 3.445 ;
        RECT  2.880 0.670 5.220 0.970 ;
        RECT  4.935 1.620 5.540 1.960 ;
        RECT  4.935 0.670 5.220 2.935 ;
        RECT  3.320 2.690 5.220 2.935 ;
    END
END XNOR2_X4_18_SVT_WB

MACRO XNOR2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.965 1.915 3.475 2.200 ;
        RECT  1.770 2.380 3.195 2.660 ;
        RECT  2.965 1.915 3.195 2.660 ;
        RECT  0.830 3.280 2.000 3.510 ;
        RECT  1.770 2.380 2.000 3.510 ;
        RECT  0.830 2.190 1.080 3.510 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.805 1.455 4.145 1.960 ;
        RECT  1.805 1.455 4.145 1.685 ;
        RECT  1.805 1.095 2.100 1.685 ;
        RECT  1.525 1.095 2.100 1.435 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.440 2.540 4.715 2.880 ;
        RECT  4.375 0.985 4.715 2.880 ;
        RECT  3.325 0.985 4.715 1.225 ;
        RECT  2.895 3.110 3.780 3.450 ;
        RECT  3.440 2.540 3.780 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.045 3.110 4.385 4.100 ;
        RECT  2.230 2.890 2.515 4.100 ;
        RECT  0.315 2.710 0.600 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.885 -0.180 2.225 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.615 0.575 0.955 1.915 ;
        RECT  0.615 1.665 1.575 1.915 ;
        RECT  1.310 1.915 2.735 2.150 ;
        RECT  1.310 1.665 1.540 3.050 ;
        RECT  2.605 0.470 4.385 0.755 ;
        RECT  2.605 0.470 2.945 1.225 ;
    END
END XNOR2_X2_18_SVT_WB

MACRO XNOR2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.180 2.970 1.540 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.810 3.760 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.660  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.965 2.380 4.330 2.720 ;
        RECT  3.990 1.225 4.330 2.720 ;
        RECT  3.200 1.225 4.330 1.455 ;
        RECT  3.200 0.870 3.540 1.455 ;
        RECT  2.440 2.955 3.250 3.295 ;
        RECT  2.965 2.380 3.250 3.295 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.960 2.990 4.300 4.100 ;
        RECT  1.680 3.015 2.020 4.100 ;
        RECT  0.200 3.005 0.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  1.680 -0.180 2.020 0.895 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.270 0.610 0.830 0.950 ;
        RECT  0.270 0.610 0.500 2.775 ;
        RECT  0.270 2.435 2.220 2.775 ;
        RECT  0.920 2.435 1.260 3.295 ;
        RECT  2.440 0.410 4.260 0.640 ;
        RECT  2.440 0.410 2.780 0.950 ;
        RECT  3.920 0.410 4.260 0.995 ;
    END
END XNOR2_X1_18_SVT_WB

MACRO XNOR2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.570 3.000 1.855 ;
        RECT  2.490 1.200 2.720 1.855 ;
        RECT  0.715 1.200 2.720 1.540 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.380 2.040 3.720 2.380 ;
        RECT  1.260 2.085 3.720 2.315 ;
        RECT  1.260 1.770 1.720 2.315 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.420 2.610 4.340 2.840 ;
        RECT  4.000 1.050 4.340 2.840 ;
        RECT  3.150 1.050 4.340 1.390 ;
        RECT  2.420 2.610 2.760 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.860 3.070 4.200 4.100 ;
        RECT  1.660 3.095 2.000 4.100 ;
        RECT  0.180 3.095 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  1.685 -0.180 2.025 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.630 0.485 2.865 ;
        RECT  0.180 2.545 2.190 2.865 ;
        RECT  0.900 2.545 1.240 3.385 ;
    END
END XNOR2_X0_18_SVT_WB

MACRO XNOR2PG_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2PG_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.210 8.925 1.735 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.553  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.770 1.455 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.375  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 3.185 7.405 3.470 ;
        RECT  5.610 0.470 7.390 0.755 ;
        RECT  0.750 0.470 7.390 0.700 ;
        RECT  0.130 0.690 4.120 0.755 ;
        RECT  0.130 2.950 2.480 3.285 ;
        RECT  0.130 0.690 0.975 0.920 ;
        RECT  0.130 0.690 0.470 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.635 2.900 11.975 4.100 ;
        RECT  10.195 3.000 10.535 4.100 ;
        RECT  8.750 3.185 9.090 4.100 ;
        RECT  1.700 3.515 2.040 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.635 -0.180 11.975 0.795 ;
        RECT  10.195 -0.180 10.535 0.740 ;
        RECT  0.180 -0.180 0.520 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  5.475 1.450 8.310 1.790 ;
        RECT  8.080 0.870 8.310 2.495 ;
        RECT  7.985 1.450 8.310 2.495 ;
        RECT  7.985 2.155 8.325 2.495 ;
        RECT  2.460 0.985 4.785 1.270 ;
        RECT  4.480 0.930 4.785 1.270 ;
        RECT  0.940 1.150 2.970 1.440 ;
        RECT  9.070 1.915 10.045 2.200 ;
        RECT  2.460 0.985 2.970 2.720 ;
        RECT  0.940 2.380 2.970 2.720 ;
        RECT  2.740 0.985 2.970 2.955 ;
        RECT  9.070 1.915 9.300 2.955 ;
        RECT  2.740 2.725 9.300 2.955 ;
        RECT  7.620 0.410 9.530 0.640 ;
        RECT  9.300 0.410 9.530 1.270 ;
        RECT  7.620 0.410 7.850 1.220 ;
        RECT  5.015 0.985 7.850 1.220 ;
        RECT  9.300 0.970 11.255 1.270 ;
        RECT  5.015 0.985 5.245 2.495 ;
        RECT  4.880 2.210 5.245 2.495 ;
        RECT  10.915 0.970 11.255 2.770 ;
        RECT  9.530 2.430 11.255 2.770 ;
    END
END XNOR2PG_X8_18_SVT_WB

MACRO XNOR2PG_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2PG_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.420 1.910 7.700 2.710 ;
        RECT  7.280 1.910 7.700 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.775 1.770 1.540 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.343  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.995 0.470 6.775 0.755 ;
        RECT  2.270 3.185 6.730 3.470 ;
        RECT  6.435 3.110 6.730 3.470 ;
        RECT  0.750 0.470 6.775 0.700 ;
        RECT  0.140 0.690 3.505 0.755 ;
        RECT  0.140 2.950 2.480 3.285 ;
        RECT  0.140 0.690 0.975 0.920 ;
        RECT  0.140 0.690 0.480 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  10.680 3.460 11.020 4.100 ;
        RECT  1.700 3.515 2.040 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  10.640 -0.180 10.980 0.810 ;
        RECT  9.200 -0.180 9.540 0.890 ;
        RECT  0.180 -0.180 0.520 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  7.780 0.880 8.215 1.680 ;
        RECT  4.860 1.450 8.215 1.680 ;
        RECT  4.860 1.450 5.145 1.790 ;
        RECT  7.930 0.880 8.215 2.940 ;
        RECT  7.195 0.410 8.805 0.650 ;
        RECT  7.195 0.410 7.535 1.220 ;
        RECT  4.400 0.985 7.535 1.220 ;
        RECT  8.480 1.120 10.260 1.440 ;
        RECT  8.480 0.410 8.805 2.720 ;
        RECT  4.400 0.985 4.630 2.495 ;
        RECT  4.265 2.210 4.630 2.495 ;
        RECT  8.480 2.380 10.260 2.720 ;
        RECT  2.460 0.985 4.170 1.270 ;
        RECT  3.865 0.930 4.170 1.270 ;
        RECT  0.940 1.150 2.970 1.440 ;
        RECT  9.035 1.810 10.830 2.150 ;
        RECT  2.460 0.985 2.970 2.720 ;
        RECT  0.940 2.380 2.970 2.720 ;
        RECT  2.740 0.985 2.970 2.955 ;
        RECT  5.715 2.615 7.190 2.880 ;
        RECT  2.740 2.725 6.055 2.955 ;
        RECT  6.960 2.615 7.190 3.510 ;
        RECT  9.925 2.950 10.830 3.230 ;
        RECT  10.490 1.810 10.830 3.230 ;
        RECT  6.960 3.170 10.265 3.510 ;
    END
END XNOR2PG_X6_18_SVT_WB

MACRO XNOR2PG_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2PG_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.575  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.470 3.675 1.760 ;
        RECT  2.940 1.080 3.280 1.760 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.820 1.120 2.250 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.350 2.230 6.285 2.515 ;
        RECT  6.055 0.700 6.285 2.515 ;
        RECT  5.350 0.700 6.285 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  1.665 3.560 2.005 4.100 ;
        RECT  0.185 2.630 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  1.665 -0.180 2.005 0.405 ;
        RECT  0.185 -0.180 0.525 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.865 1.005 4.245 1.290 ;
        RECT  3.970 1.520 5.825 1.860 ;
        RECT  3.970 1.005 4.245 2.515 ;
        RECT  3.905 2.230 4.245 2.515 ;
        RECT  2.425 0.470 4.970 0.775 ;
        RECT  2.425 0.470 2.700 2.815 ;
        RECT  2.425 2.475 2.935 2.815 ;
        RECT  2.705 2.745 6.410 2.975 ;
        RECT  0.905 0.590 1.245 1.345 ;
        RECT  0.905 1.115 2.100 1.345 ;
        RECT  6.515 0.480 6.800 2.515 ;
        RECT  1.815 1.115 2.100 3.330 ;
        RECT  0.905 2.630 2.100 3.330 ;
        RECT  0.905 3.045 2.485 3.330 ;
        RECT  6.745 2.175 7.085 3.510 ;
        RECT  2.235 3.205 7.085 3.510 ;
    END
END XNOR2PG_X4_18_SVT_WB

MACRO XNOR2PG_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2PG_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.602  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.260 2.710 1.810 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.200 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 2.230 5.385 2.515 ;
        RECT  5.155 0.700 5.385 2.515 ;
        RECT  4.450 0.700 5.385 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  0.940 3.460 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  0.940 -0.180 1.280 0.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.005 1.520 4.925 1.860 ;
        RECT  3.005 1.005 3.370 2.515 ;
        RECT  1.700 0.470 4.070 0.775 ;
        RECT  1.700 0.470 1.940 2.760 ;
        RECT  1.700 2.450 2.210 2.760 ;
        RECT  1.980 2.745 5.510 2.975 ;
        RECT  0.180 0.535 0.520 1.460 ;
        RECT  0.180 1.230 1.470 1.460 ;
        RECT  5.615 0.480 5.900 2.015 ;
        RECT  0.180 2.575 1.470 2.915 ;
        RECT  1.160 1.230 1.470 3.230 ;
        RECT  1.160 2.990 1.750 3.230 ;
        RECT  0.180 2.575 0.520 3.275 ;
        RECT  5.740 1.690 6.045 3.490 ;
        RECT  1.510 3.205 6.045 3.490 ;
    END
END XNOR2PG_X2_18_SVT_WB

MACRO XNOR2PG_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN XNOR2PG_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.602  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.260 2.710 1.810 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.200 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 2.230 5.385 2.515 ;
        RECT  5.155 0.700 5.385 2.515 ;
        RECT  4.450 0.700 5.385 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  0.940 3.460 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  0.940 -0.180 1.280 0.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.005 1.520 4.925 1.860 ;
        RECT  3.005 1.005 3.370 2.515 ;
        RECT  1.700 0.470 4.070 0.775 ;
        RECT  1.700 0.470 1.940 2.760 ;
        RECT  1.700 2.450 2.210 2.760 ;
        RECT  1.980 2.745 5.510 2.975 ;
        RECT  0.180 0.535 0.520 1.460 ;
        RECT  0.180 1.230 1.470 1.460 ;
        RECT  5.615 0.480 5.900 2.015 ;
        RECT  0.180 2.575 1.470 2.915 ;
        RECT  1.160 1.230 1.470 3.230 ;
        RECT  1.160 2.990 1.750 3.230 ;
        RECT  5.740 1.690 6.045 3.490 ;
        RECT  1.510 3.205 6.045 3.490 ;
    END
END XNOR2PG_X1_18_SVT_WB

MACRO TLAT_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLAT_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.080 1.810 1.590 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.327  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.110 2.775 2.555 ;
        RECT  0.690 2.095 2.775 2.325 ;
        RECT  2.190 1.110 2.775 2.325 ;
        RECT  0.690 1.155 1.030 2.325 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.740 1.100 6.080 2.720 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.195 0.470 7.700 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.930 2.640 8.220 4.100 ;
        RECT  3.640 3.000 3.980 4.100 ;
        RECT  0.940 3.515 1.660 4.100 ;
        RECT  0.940 3.185 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.930 -0.180 8.220 1.280 ;
        RECT  3.640 -0.180 3.980 0.810 ;
        RECT  1.220 -0.180 1.560 0.850 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.570 0.800 0.910 ;
        RECT  0.180 0.570 0.460 2.955 ;
        RECT  0.180 2.615 2.230 2.955 ;
        RECT  1.890 2.615 2.230 3.475 ;
        RECT  2.410 0.570 3.235 0.880 ;
        RECT  3.005 1.455 5.400 1.685 ;
        RECT  4.120 1.455 5.400 1.960 ;
        RECT  3.005 0.570 3.235 3.275 ;
        RECT  2.460 2.935 3.235 3.275 ;
        RECT  4.360 0.525 6.965 0.865 ;
        RECT  4.360 0.525 4.700 1.225 ;
        RECT  3.465 1.915 3.790 2.495 ;
        RECT  3.465 2.265 4.700 2.495 ;
        RECT  4.360 2.265 4.700 3.245 ;
        RECT  6.680 0.525 6.965 3.245 ;
        RECT  4.360 2.950 6.965 3.245 ;
    END
END TLAT_X4_18_SVT_WB

MACRO TLAT_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLAT_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.070 1.660 1.540 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.327  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.065 1.120 2.545 2.510 ;
        RECT  0.575 1.820 2.545 2.110 ;
        RECT  2.040 1.120 2.545 2.110 ;
        RECT  0.575 1.225 0.860 2.110 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.845 2.375 5.460 2.760 ;
        RECT  5.155 1.020 5.460 2.760 ;
        RECT  4.845 1.020 5.460 1.395 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.245 0.470 6.580 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  3.330 3.495 3.670 4.100 ;
        RECT  0.940 3.445 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  1.040 -0.180 1.380 0.835 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.550 0.620 0.890 ;
        RECT  0.115 0.550 0.345 3.165 ;
        RECT  0.115 2.705 0.520 3.165 ;
        RECT  0.115 2.935 2.050 3.165 ;
        RECT  1.710 2.935 2.050 3.510 ;
        RECT  2.230 0.550 3.005 0.890 ;
        RECT  2.775 1.240 4.615 1.580 ;
        RECT  4.310 1.240 4.615 2.000 ;
        RECT  2.775 0.550 3.005 3.365 ;
        RECT  2.280 3.025 3.005 3.365 ;
        RECT  4.090 0.550 6.015 0.790 ;
        RECT  4.090 0.550 4.430 0.890 ;
        RECT  3.235 1.880 3.520 2.860 ;
        RECT  3.235 2.630 4.150 2.860 ;
        RECT  3.920 2.630 4.150 3.330 ;
        RECT  5.720 0.550 6.015 3.330 ;
        RECT  3.920 2.990 6.015 3.330 ;
    END
END TLAT_X2_18_SVT_WB

MACRO TLAT_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLAT_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.090 1.590 1.540 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.327  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.985 2.170 2.575 2.695 ;
        RECT  2.290 1.135 2.575 2.695 ;
        RECT  1.820 1.135 2.575 1.590 ;
        RECT  0.575 2.170 2.575 2.400 ;
        RECT  0.575 1.590 0.890 2.400 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.875 1.080 5.215 2.820 ;
        RECT  4.620 1.080 5.215 1.590 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 2.650 6.580 3.095 ;
        RECT  6.300 1.005 6.580 3.095 ;
        RECT  6.200 1.005 6.580 1.345 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  5.635 3.525 6.445 4.100 ;
        RECT  0.990 3.445 1.330 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  5.635 -0.180 6.445 0.380 ;
        RECT  1.115 -0.180 1.455 0.855 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.570 0.655 0.910 ;
        RECT  0.115 0.570 0.345 3.165 ;
        RECT  0.115 2.705 0.520 3.165 ;
        RECT  0.115 2.935 2.060 3.165 ;
        RECT  1.720 2.935 2.060 3.510 ;
        RECT  2.265 0.570 3.035 0.905 ;
        RECT  2.805 1.245 4.295 1.545 ;
        RECT  3.955 1.245 4.295 2.000 ;
        RECT  2.805 0.570 3.035 3.155 ;
        RECT  2.290 2.925 3.035 3.155 ;
        RECT  2.290 2.925 2.580 3.435 ;
        RECT  4.175 0.610 5.845 0.850 ;
        RECT  5.615 1.545 6.070 2.355 ;
        RECT  3.265 1.775 3.605 2.700 ;
        RECT  3.265 2.470 4.235 2.700 ;
        RECT  4.005 2.470 4.235 3.295 ;
        RECT  5.615 0.610 5.845 3.295 ;
        RECT  4.005 3.050 5.845 3.295 ;
    END
END TLAT_X1_18_SVT_WB

MACRO TLATSR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATSR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.820 3.270 2.100 ;
        RECT  2.520 1.820 2.860 2.250 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.291  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.905 1.350 4.135 2.730 ;
        RECT  1.180 1.350 4.135 1.580 ;
        RECT  2.890 1.260 3.270 1.580 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.220 2.330 10.860 3.295 ;
        RECT  10.630 0.575 10.860 3.295 ;
        RECT  10.575 0.575 10.860 1.445 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.930 2.380 9.340 2.705 ;
        RECT  9.000 0.630 9.340 2.705 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.810 2.210 2.270 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.690 2.105 6.245 2.660 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  11.215 2.375 11.600 4.100 ;
        RECT  9.730 3.570 10.145 4.100 ;
        RECT  6.395 3.570 6.735 4.100 ;
        RECT  4.935 2.965 5.165 4.100 ;
        RECT  0.995 3.515 1.225 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  11.210 -0.180 11.615 1.470 ;
        RECT  9.815 -0.180 10.045 0.875 ;
        RECT  5.105 -0.180 5.335 1.240 ;
        RECT  1.565 -0.180 1.795 1.035 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.235 0.775 0.905 1.115 ;
        RECT  3.180 2.400 3.535 2.735 ;
        RECT  0.235 2.505 3.535 2.735 ;
        RECT  0.235 0.775 0.465 3.430 ;
        RECT  3.445 0.705 4.595 1.045 ;
        RECT  4.365 2.335 5.440 2.675 ;
        RECT  4.365 0.705 4.595 3.305 ;
        RECT  1.665 2.965 4.595 3.305 ;
        RECT  4.825 1.645 6.685 1.875 ;
        RECT  6.255 0.980 6.685 1.875 ;
        RECT  4.825 1.645 5.055 2.005 ;
        RECT  6.475 1.780 7.210 2.120 ;
        RECT  6.475 1.780 6.705 3.285 ;
        RECT  5.690 2.945 6.705 3.285 ;
        RECT  7.470 1.100 7.940 1.440 ;
        RECT  9.670 1.740 10.400 2.085 ;
        RECT  7.470 1.100 7.700 3.285 ;
        RECT  7.210 2.845 7.700 3.285 ;
        RECT  9.670 1.740 9.900 3.285 ;
        RECT  7.210 3.035 9.900 3.285 ;
    END
END TLATSR_X4_18_SVT_WB

MACRO TLATSR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATSR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.820 3.270 2.100 ;
        RECT  2.520 1.820 2.860 2.250 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.291  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.905 1.350 4.135 2.730 ;
        RECT  1.180 1.350 4.135 1.580 ;
        RECT  2.890 1.260 3.270 1.580 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.610 2.365 10.195 3.295 ;
        RECT  9.965 0.575 10.195 3.295 ;
        RECT  9.910 0.575 10.195 1.445 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.930 2.380 8.675 2.705 ;
        RECT  8.335 0.630 8.675 2.705 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.810 2.210 2.270 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.690 2.105 6.245 2.660 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.065 3.570 9.480 4.100 ;
        RECT  6.395 3.570 6.735 4.100 ;
        RECT  4.935 2.965 5.165 4.100 ;
        RECT  0.995 3.515 1.225 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.150 -0.180 9.380 0.875 ;
        RECT  5.105 -0.180 5.335 1.240 ;
        RECT  1.565 -0.180 1.795 1.035 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.235 0.775 0.905 1.115 ;
        RECT  3.185 2.400 3.530 2.735 ;
        RECT  0.235 2.505 3.530 2.735 ;
        RECT  0.235 0.775 0.465 3.430 ;
        RECT  3.445 0.705 4.595 1.045 ;
        RECT  4.365 2.335 5.440 2.675 ;
        RECT  4.365 0.705 4.595 3.305 ;
        RECT  1.665 2.965 4.595 3.305 ;
        RECT  4.825 1.645 6.685 1.875 ;
        RECT  6.255 0.980 6.685 1.875 ;
        RECT  4.825 1.645 5.055 2.005 ;
        RECT  6.475 1.780 7.210 2.120 ;
        RECT  6.475 1.780 6.705 3.285 ;
        RECT  5.690 2.945 6.705 3.285 ;
        RECT  7.470 1.100 7.940 1.440 ;
        RECT  9.080 1.740 9.735 2.130 ;
        RECT  7.470 1.100 7.700 3.285 ;
        RECT  7.210 2.845 7.700 3.285 ;
        RECT  9.080 1.740 9.370 3.285 ;
        RECT  7.210 3.035 9.370 3.285 ;
    END
END TLATSR_X2_18_SVT_WB

MACRO TLATSR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATSR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.820 3.270 2.100 ;
        RECT  2.520 1.820 2.860 2.250 ;
        END
    END D
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.291  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.905 1.350 4.135 2.730 ;
        RECT  1.180 1.350 4.135 1.580 ;
        RECT  2.890 1.260 3.270 1.580 ;
        END
    END G
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.610 2.365 10.195 2.665 ;
        RECT  9.965 0.575 10.195 2.665 ;
        RECT  9.910 0.575 10.195 0.915 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.930 2.380 8.675 2.705 ;
        RECT  8.335 0.630 8.675 2.705 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.810 2.210 2.270 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.690 2.105 6.245 2.660 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.065 3.570 9.480 4.100 ;
        RECT  6.395 3.570 6.735 4.100 ;
        RECT  4.935 2.965 5.165 4.100 ;
        RECT  0.995 3.515 1.225 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.150 -0.180 9.380 0.875 ;
        RECT  5.105 -0.180 5.335 1.240 ;
        RECT  1.565 -0.180 1.795 1.035 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.235 0.775 0.905 1.115 ;
        RECT  3.195 2.400 3.530 2.735 ;
        RECT  0.235 2.505 3.530 2.735 ;
        RECT  0.235 0.775 0.465 3.430 ;
        RECT  3.445 0.705 4.595 1.045 ;
        RECT  4.365 2.335 5.440 2.675 ;
        RECT  4.365 0.705 4.595 3.305 ;
        RECT  1.665 2.965 4.595 3.305 ;
        RECT  4.825 1.645 6.685 1.875 ;
        RECT  6.255 0.980 6.685 1.875 ;
        RECT  4.825 1.645 5.055 2.005 ;
        RECT  6.475 1.780 7.210 2.120 ;
        RECT  6.475 1.780 6.705 3.285 ;
        RECT  5.690 2.945 6.705 3.285 ;
        RECT  7.470 1.100 7.940 1.440 ;
        RECT  9.080 1.105 9.735 1.495 ;
        RECT  7.470 1.100 7.700 3.285 ;
        RECT  7.210 2.845 7.700 3.285 ;
        RECT  9.080 1.105 9.370 3.285 ;
        RECT  7.210 3.035 9.370 3.285 ;
    END
END TLATSR_X1_18_SVT_WB

MACRO TLATN_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATN_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.105 1.775 1.590 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.287  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.890 2.750 2.180 3.480 ;
        RECT  1.105 2.750 2.180 2.980 ;
        RECT  1.105 2.025 1.360 2.980 ;
        RECT  0.690 2.025 1.360 2.365 ;
        RECT  0.690 1.195 1.030 2.365 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.740 1.100 6.080 2.720 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.195 0.470 7.700 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.930 2.640 8.220 4.100 ;
        RECT  3.710 3.420 4.050 4.100 ;
        RECT  0.945 3.515 1.660 4.100 ;
        RECT  0.945 3.210 1.285 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.930 -0.180 8.220 1.280 ;
        RECT  3.710 -0.180 4.050 0.410 ;
        RECT  1.220 -0.180 1.560 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.185 0.635 2.235 0.875 ;
        RECT  2.005 0.635 2.235 1.470 ;
        RECT  2.005 1.160 2.835 1.470 ;
        RECT  2.495 1.160 2.835 2.535 ;
        RECT  0.185 0.635 0.460 2.955 ;
        RECT  0.185 2.615 0.525 2.955 ;
        RECT  2.465 0.590 3.295 0.930 ;
        RECT  3.065 1.475 5.455 1.705 ;
        RECT  4.285 1.475 5.455 1.960 ;
        RECT  3.065 0.590 3.295 2.995 ;
        RECT  2.415 2.765 3.295 2.995 ;
        RECT  2.415 2.765 2.755 3.275 ;
        RECT  4.470 0.530 6.965 0.870 ;
        RECT  4.470 0.530 4.810 1.245 ;
        RECT  3.560 1.935 3.900 2.460 ;
        RECT  3.560 2.230 4.810 2.460 ;
        RECT  4.470 2.230 4.810 3.210 ;
        RECT  6.680 0.530 6.965 3.210 ;
        RECT  4.470 2.950 6.965 3.210 ;
    END
END TLATN_X4_18_SVT_WB

MACRO TLATN_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATN_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.165 1.070 1.595 1.540 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.285  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.510 3.225 2.180 3.510 ;
        RECT  1.210 2.030 1.845 3.225 ;
        RECT  0.575 2.030 1.845 2.370 ;
        RECT  0.575 1.090 0.860 2.370 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.850 2.300 5.460 2.720 ;
        RECT  5.100 1.100 5.460 2.720 ;
        RECT  4.850 1.100 5.460 1.445 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.225 0.470 6.580 3.450 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  3.340 3.405 3.680 4.100 ;
        RECT  0.940 3.455 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  1.040 -0.180 1.380 0.380 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.535 0.620 0.840 ;
        RECT  0.115 0.610 2.055 0.840 ;
        RECT  1.825 0.610 2.055 1.410 ;
        RECT  1.825 1.105 2.555 1.410 ;
        RECT  2.265 1.105 2.555 2.510 ;
        RECT  0.115 0.535 0.345 3.155 ;
        RECT  0.115 2.815 0.520 3.155 ;
        RECT  2.285 0.535 3.015 0.875 ;
        RECT  2.785 1.230 4.155 1.470 ;
        RECT  3.860 1.230 4.155 1.980 ;
        RECT  3.860 1.640 4.620 1.980 ;
        RECT  2.785 0.535 3.015 2.990 ;
        RECT  2.190 2.740 3.015 2.990 ;
        RECT  4.100 0.550 5.995 0.790 ;
        RECT  4.100 0.550 4.440 0.890 ;
        RECT  3.245 2.150 3.530 2.680 ;
        RECT  3.245 2.450 4.440 2.680 ;
        RECT  4.095 2.450 4.440 3.190 ;
        RECT  5.710 0.550 5.995 3.190 ;
        RECT  4.095 2.950 5.995 3.190 ;
    END
END TLATN_X2_18_SVT_WB

MACRO TLATN_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATN_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.090 1.570 1.660 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.287  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.690 2.935 2.030 3.510 ;
        RECT  1.240 2.935 2.030 3.165 ;
        RECT  1.240 2.170 1.555 3.165 ;
        RECT  0.575 2.170 1.555 2.400 ;
        RECT  0.575 1.590 0.890 2.400 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.875 1.080 5.215 2.820 ;
        RECT  4.620 1.080 5.215 1.590 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 2.650 6.580 3.095 ;
        RECT  6.300 1.005 6.580 3.095 ;
        RECT  6.200 1.005 6.580 1.345 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  5.635 3.515 6.445 4.100 ;
        RECT  0.940 3.430 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  5.635 -0.180 6.445 0.350 ;
        RECT  0.955 -0.180 1.360 0.365 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.615 2.030 0.855 ;
        RECT  1.800 0.615 2.030 1.475 ;
        RECT  1.800 1.175 2.575 1.475 ;
        RECT  0.115 0.615 0.345 3.165 ;
        RECT  2.290 1.175 2.575 2.695 ;
        RECT  0.115 2.690 0.520 3.165 ;
        RECT  2.260 0.540 3.035 0.945 ;
        RECT  2.805 1.165 4.390 1.505 ;
        RECT  4.050 1.165 4.390 1.975 ;
        RECT  2.805 0.540 3.035 3.155 ;
        RECT  2.260 2.925 3.035 3.155 ;
        RECT  2.260 2.925 2.550 3.435 ;
        RECT  4.175 0.580 5.845 0.850 ;
        RECT  5.615 1.545 6.070 2.355 ;
        RECT  3.265 1.870 3.605 2.850 ;
        RECT  3.265 2.620 4.515 2.850 ;
        RECT  5.615 0.580 5.845 3.280 ;
        RECT  4.175 3.050 5.845 3.280 ;
        RECT  4.175 2.620 4.515 3.435 ;
    END
END TLATN_X1_18_SVT_WB

MACRO TLATNTSCA_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.480  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.015 1.680 7.795 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.705 1.610 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.800 1.725 11.205 3.410 ;
        RECT  10.830 0.540 11.205 3.410 ;
        RECT  9.430 1.725 11.205 2.175 ;
        RECT  9.430 1.725 9.805 3.445 ;
        RECT  9.430 0.490 9.780 3.445 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.500 0.980 2.405 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.560 2.615 11.900 4.100 ;
        RECT  10.170 2.635 10.460 4.100 ;
        RECT  6.010 3.440 6.820 4.100 ;
        RECT  3.580 2.690 3.920 4.100 ;
        RECT  0.190 2.640 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.560 -0.180 11.900 1.385 ;
        RECT  10.170 -0.180 10.460 1.300 ;
        RECT  5.760 -0.180 6.100 0.410 ;
        RECT  3.580 -0.180 3.920 1.375 ;
        RECT  1.005 -0.180 1.705 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.645 0.530 1.005 ;
        RECT  0.190 0.775 1.795 1.005 ;
        RECT  1.510 0.775 1.795 1.405 ;
        RECT  2.025 0.545 2.255 3.510 ;
        RECT  2.025 3.210 2.960 3.510 ;
        RECT  2.485 2.120 4.345 2.460 ;
        RECT  2.485 1.085 2.770 2.980 ;
        RECT  4.810 0.490 5.320 0.835 ;
        RECT  5.035 0.490 5.320 2.950 ;
        RECT  5.570 1.650 6.765 1.990 ;
        RECT  6.480 1.085 6.765 2.750 ;
        RECT  4.300 1.085 4.640 1.890 ;
        RECT  3.360 1.605 4.805 1.890 ;
        RECT  8.220 1.695 8.585 2.690 ;
        RECT  6.995 2.460 8.585 2.690 ;
        RECT  4.575 1.555 4.805 3.410 ;
        RECT  4.300 2.690 4.805 3.410 ;
        RECT  5.550 2.980 7.225 3.210 ;
        RECT  6.995 2.460 7.225 3.210 ;
        RECT  4.300 3.180 5.780 3.410 ;
        RECT  7.180 0.515 7.520 1.355 ;
        RECT  7.180 1.100 9.200 1.355 ;
        RECT  8.915 1.100 9.200 3.445 ;
        RECT  8.050 3.105 9.200 3.445 ;
    END
END TLATNTSCA_X8_18_SVT_WB

MACRO TLATNTSCA_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.480  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.995 1.680 7.730 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.705 1.610 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.239  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.890 2.480 11.235 3.445 ;
        RECT  9.430 1.125 11.235 1.360 ;
        RECT  10.890 0.490 11.235 1.360 ;
        RECT  9.430 2.480 11.235 2.740 ;
        RECT  10.215 1.125 10.660 2.740 ;
        RECT  9.430 2.480 9.810 3.460 ;
        RECT  9.430 0.490 9.805 1.360 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.500 0.980 2.405 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  10.200 3.045 10.510 4.100 ;
        RECT  6.010 3.440 6.820 4.100 ;
        RECT  3.580 2.690 3.920 4.100 ;
        RECT  0.190 2.640 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  10.160 -0.180 10.500 0.845 ;
        RECT  5.760 -0.180 6.100 0.410 ;
        RECT  3.580 -0.180 3.920 1.375 ;
        RECT  1.005 -0.180 1.705 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.645 0.530 1.005 ;
        RECT  0.190 0.775 1.795 1.005 ;
        RECT  1.510 0.775 1.795 1.405 ;
        RECT  2.025 0.545 2.255 3.510 ;
        RECT  2.025 3.210 2.960 3.510 ;
        RECT  2.485 2.120 4.345 2.460 ;
        RECT  2.485 1.085 2.770 2.980 ;
        RECT  4.810 0.490 5.320 0.835 ;
        RECT  5.035 0.490 5.320 2.950 ;
        RECT  5.570 1.650 6.765 1.990 ;
        RECT  6.480 1.085 6.765 2.750 ;
        RECT  4.300 1.085 4.640 1.890 ;
        RECT  3.360 1.605 4.805 1.890 ;
        RECT  8.245 1.755 8.585 2.690 ;
        RECT  6.995 2.460 8.585 2.690 ;
        RECT  4.575 1.555 4.805 3.410 ;
        RECT  4.300 2.690 4.805 3.410 ;
        RECT  5.550 2.980 7.225 3.210 ;
        RECT  6.995 2.460 7.225 3.210 ;
        RECT  4.300 3.180 5.780 3.410 ;
        RECT  7.180 0.565 7.535 1.380 ;
        RECT  7.180 1.110 9.200 1.380 ;
        RECT  8.950 1.670 9.735 1.910 ;
        RECT  8.950 1.110 9.200 3.445 ;
        RECT  8.050 3.105 9.200 3.445 ;
    END
END TLATNTSCA_X6_18_SVT_WB

MACRO TLATNTSCA_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.065 1.210 7.700 1.760 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.705 1.610 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.870 0.490 9.380 3.445 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.500 0.980 2.405 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  9.610 2.635 9.900 4.100 ;
        RECT  6.010 3.440 6.820 4.100 ;
        RECT  3.580 2.690 3.920 4.100 ;
        RECT  0.190 2.640 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  9.610 -0.180 9.900 1.300 ;
        RECT  5.760 -0.180 6.100 0.820 ;
        RECT  3.580 -0.180 3.920 1.375 ;
        RECT  1.005 -0.180 1.705 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.645 0.530 1.005 ;
        RECT  0.190 0.775 1.795 1.005 ;
        RECT  1.510 0.775 1.795 1.405 ;
        RECT  2.025 0.545 2.255 3.510 ;
        RECT  2.025 3.210 2.960 3.510 ;
        RECT  2.485 2.120 4.345 2.460 ;
        RECT  2.485 1.085 2.770 2.980 ;
        RECT  4.810 0.560 5.320 0.900 ;
        RECT  5.035 0.560 5.320 2.950 ;
        RECT  5.570 1.650 6.765 1.990 ;
        RECT  6.480 1.130 6.765 2.750 ;
        RECT  4.300 1.085 4.640 1.890 ;
        RECT  3.360 1.605 4.805 1.890 ;
        RECT  7.640 2.095 7.980 2.875 ;
        RECT  6.995 2.535 7.980 2.875 ;
        RECT  4.575 1.555 4.805 3.410 ;
        RECT  4.300 2.690 4.805 3.410 ;
        RECT  5.550 2.980 7.225 3.210 ;
        RECT  6.995 2.535 7.225 3.210 ;
        RECT  4.300 3.180 5.780 3.410 ;
        RECT  6.560 0.430 8.640 0.770 ;
        RECT  8.355 0.430 8.640 3.445 ;
        RECT  7.455 3.105 8.640 3.445 ;
    END
END TLATNTSCA_X4_18_SVT_WB

MACRO TLATNTSCA_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.065 1.210 7.700 1.760 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.705 1.610 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.894  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.870 0.490 9.380 3.445 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.500 0.980 2.405 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  9.610 2.785 9.900 4.100 ;
        RECT  6.010 3.440 6.820 4.100 ;
        RECT  3.580 2.690 3.920 4.100 ;
        RECT  0.190 2.640 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  9.610 -0.180 9.900 0.960 ;
        RECT  5.760 -0.180 6.100 0.820 ;
        RECT  3.580 -0.180 3.920 1.375 ;
        RECT  1.005 -0.180 1.705 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.645 0.530 1.005 ;
        RECT  0.190 0.775 1.795 1.005 ;
        RECT  1.510 0.775 1.795 1.405 ;
        RECT  2.025 0.545 2.255 3.510 ;
        RECT  2.025 3.210 2.960 3.510 ;
        RECT  2.485 2.120 4.345 2.460 ;
        RECT  2.485 1.085 2.770 2.980 ;
        RECT  4.810 0.560 5.320 0.900 ;
        RECT  5.035 0.560 5.320 2.950 ;
        RECT  5.570 1.650 6.765 1.990 ;
        RECT  6.480 1.130 6.765 2.750 ;
        RECT  4.300 1.085 4.640 1.890 ;
        RECT  3.360 1.605 4.805 1.890 ;
        RECT  7.640 2.095 7.980 2.875 ;
        RECT  6.995 2.535 7.980 2.875 ;
        RECT  4.575 1.555 4.805 3.410 ;
        RECT  4.300 2.690 4.805 3.410 ;
        RECT  5.550 2.980 7.225 3.210 ;
        RECT  6.995 2.535 7.225 3.210 ;
        RECT  4.300 3.180 5.780 3.410 ;
        RECT  6.560 0.430 8.640 0.770 ;
        RECT  8.355 0.430 8.640 3.445 ;
        RECT  7.455 3.105 8.640 3.445 ;
    END
END TLATNTSCA_X3_18_SVT_WB

MACRO TLATNTSCA_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.160 1.105 8.030 1.860 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.565 1.710 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.054  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.870 0.470 9.380 3.460 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.197  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.450 0.710 2.260 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  6.280 3.545 6.735 4.100 ;
        RECT  3.610 2.605 3.950 4.100 ;
        RECT  0.210 2.555 0.550 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  8.110 -0.180 8.450 0.415 ;
        RECT  5.815 -0.180 6.155 0.900 ;
        RECT  3.610 -0.180 3.950 1.290 ;
        RECT  0.970 -0.180 1.725 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.210 0.560 0.550 1.020 ;
        RECT  0.210 0.790 1.825 1.020 ;
        RECT  1.540 0.790 1.825 1.320 ;
        RECT  2.055 0.460 2.285 3.510 ;
        RECT  2.055 3.170 3.025 3.510 ;
        RECT  2.515 2.035 4.375 2.375 ;
        RECT  2.515 1.000 2.800 2.895 ;
        RECT  4.840 0.505 5.370 0.825 ;
        RECT  5.065 0.505 5.370 2.970 ;
        RECT  5.600 1.805 6.795 2.315 ;
        RECT  6.510 1.130 6.795 2.750 ;
        RECT  4.330 1.055 4.835 1.805 ;
        RECT  3.390 1.520 4.835 1.805 ;
        RECT  7.025 2.440 7.990 2.775 ;
        RECT  4.605 1.055 4.835 3.430 ;
        RECT  4.330 2.605 4.835 3.430 ;
        RECT  5.665 3.085 7.255 3.315 ;
        RECT  7.025 2.440 7.255 3.315 ;
        RECT  4.330 3.200 5.910 3.430 ;
        RECT  6.640 0.430 6.980 0.875 ;
        RECT  6.640 0.645 8.600 0.875 ;
        RECT  8.260 0.645 8.600 3.445 ;
        RECT  7.485 3.105 8.600 3.445 ;
    END
END TLATNTSCA_X2_18_SVT_WB

MACRO TLATNTSCA_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.080 1.680 9.295 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.075 1.705 1.610 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.926  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.770 0.490 18.110 3.355 ;
        RECT  12.280 1.725 18.110 2.170 ;
        RECT  16.450 0.555 16.790 3.355 ;
        RECT  15.010 0.570 15.350 3.410 ;
        RECT  13.650 1.725 14.055 3.410 ;
        RECT  13.680 0.540 14.055 3.410 ;
        RECT  12.280 1.725 14.055 2.175 ;
        RECT  12.280 1.725 12.660 3.445 ;
        RECT  12.280 0.490 12.650 3.445 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.500 0.785 2.405 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 19.040 4.100 ;
        RECT  18.490 2.565 18.830 4.100 ;
        RECT  15.730 2.495 16.070 4.100 ;
        RECT  12.970 2.635 13.310 4.100 ;
        RECT  6.075 3.440 7.415 4.100 ;
        RECT  3.580 2.690 3.920 4.100 ;
        RECT  0.190 2.640 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 19.040 0.180 ;
        RECT  18.490 -0.180 18.830 1.270 ;
        RECT  15.730 -0.180 16.070 1.285 ;
        RECT  12.970 -0.180 13.310 1.300 ;
        RECT  5.825 -0.180 6.165 0.415 ;
        RECT  3.645 -0.180 3.985 1.185 ;
        RECT  1.005 -0.180 1.705 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.645 0.530 1.005 ;
        RECT  0.190 0.775 1.795 1.005 ;
        RECT  1.510 0.775 1.795 1.405 ;
        RECT  2.025 0.545 2.255 3.510 ;
        RECT  2.025 3.210 2.960 3.510 ;
        RECT  4.180 1.875 4.410 2.460 ;
        RECT  2.485 2.120 4.410 2.460 ;
        RECT  2.485 1.085 2.770 2.980 ;
        RECT  4.875 0.430 5.385 0.770 ;
        RECT  5.100 0.430 5.385 2.950 ;
        RECT  5.635 1.650 6.830 1.990 ;
        RECT  6.545 1.070 6.830 2.750 ;
        RECT  7.955 0.540 11.190 0.820 ;
        RECT  4.365 1.085 4.870 1.645 ;
        RECT  3.360 1.415 4.870 1.645 ;
        RECT  3.360 1.415 3.705 1.890 ;
        RECT  9.905 1.710 11.235 2.040 ;
        RECT  9.905 1.710 10.245 2.770 ;
        RECT  7.275 2.535 10.245 2.770 ;
        RECT  4.640 1.085 4.870 3.410 ;
        RECT  4.365 2.690 4.870 3.410 ;
        RECT  5.615 2.980 7.505 3.210 ;
        RECT  7.275 2.535 7.505 3.210 ;
        RECT  4.365 3.180 5.845 3.410 ;
        RECT  7.245 0.515 7.585 1.355 ;
        RECT  7.245 1.100 12.050 1.355 ;
        RECT  11.765 1.100 12.050 3.255 ;
        RECT  7.960 3.025 12.050 3.255 ;
    END
END TLATNTSCA_X20_18_SVT_WB

MACRO TLATNTSCA_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.080 1.680 9.295 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.705 1.610 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.741  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.450 0.555 16.790 3.355 ;
        RECT  12.280 1.725 16.790 2.170 ;
        RECT  15.010 0.570 15.350 3.410 ;
        RECT  13.650 1.725 14.055 3.410 ;
        RECT  13.680 0.540 14.055 3.410 ;
        RECT  12.280 1.725 14.055 2.175 ;
        RECT  12.280 1.725 12.660 3.445 ;
        RECT  12.280 0.490 12.650 3.445 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.500 0.790 2.405 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  17.170 2.540 17.510 4.100 ;
        RECT  15.730 2.495 16.070 4.100 ;
        RECT  12.970 2.635 13.310 4.100 ;
        RECT  6.075 3.440 7.415 4.100 ;
        RECT  3.580 2.690 3.920 4.100 ;
        RECT  0.190 2.640 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  17.170 -0.180 17.510 1.325 ;
        RECT  15.730 -0.180 16.070 1.285 ;
        RECT  12.970 -0.180 13.310 1.300 ;
        RECT  5.825 -0.180 6.165 0.415 ;
        RECT  3.645 -0.180 3.985 1.185 ;
        RECT  1.005 -0.180 1.705 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.645 0.530 1.005 ;
        RECT  0.190 0.775 1.795 1.005 ;
        RECT  1.510 0.775 1.795 1.405 ;
        RECT  2.025 0.545 2.255 3.510 ;
        RECT  2.025 3.210 2.960 3.510 ;
        RECT  4.180 1.875 4.410 2.460 ;
        RECT  2.485 2.120 4.410 2.460 ;
        RECT  2.485 1.085 2.770 2.980 ;
        RECT  4.875 0.430 5.385 0.770 ;
        RECT  5.100 0.430 5.385 2.950 ;
        RECT  5.635 1.650 6.830 1.990 ;
        RECT  6.545 1.070 6.830 2.750 ;
        RECT  7.955 0.540 11.190 0.820 ;
        RECT  4.365 1.085 4.870 1.645 ;
        RECT  3.360 1.415 4.870 1.645 ;
        RECT  3.360 1.415 3.705 1.890 ;
        RECT  9.905 1.710 11.235 2.040 ;
        RECT  9.905 1.710 10.245 2.770 ;
        RECT  7.275 2.535 10.245 2.770 ;
        RECT  4.640 1.085 4.870 3.410 ;
        RECT  4.365 2.690 4.870 3.410 ;
        RECT  5.615 2.980 7.505 3.210 ;
        RECT  7.275 2.535 7.505 3.210 ;
        RECT  4.365 3.180 5.845 3.410 ;
        RECT  7.245 0.515 7.585 1.355 ;
        RECT  7.245 1.100 12.050 1.355 ;
        RECT  11.765 1.100 12.050 3.255 ;
        RECT  7.960 3.025 12.050 3.255 ;
    END
END TLATNTSCA_X16_18_SVT_WB

MACRO TLATNTSCA_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNTSCA_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.080 1.680 9.295 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.705 1.610 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.556  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.130 0.570 15.470 3.410 ;
        RECT  12.280 1.725 15.470 2.170 ;
        RECT  13.650 1.725 14.055 3.410 ;
        RECT  13.680 0.540 14.055 3.410 ;
        RECT  12.280 1.725 14.055 2.175 ;
        RECT  12.280 1.725 12.660 3.445 ;
        RECT  12.280 0.490 12.650 3.445 ;
        END
    END ECK
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.500 0.775 2.405 ;
        END
    END SE
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  14.410 2.600 14.750 4.100 ;
        RECT  12.970 2.635 13.310 4.100 ;
        RECT  6.075 3.440 7.415 4.100 ;
        RECT  3.580 2.690 3.920 4.100 ;
        RECT  0.190 2.640 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  14.410 -0.180 14.750 1.295 ;
        RECT  12.970 -0.180 13.310 1.300 ;
        RECT  5.825 -0.180 6.165 0.415 ;
        RECT  3.645 -0.180 3.985 1.185 ;
        RECT  1.005 -0.180 1.705 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.645 0.530 1.005 ;
        RECT  0.190 0.775 1.795 1.005 ;
        RECT  1.510 0.775 1.795 1.405 ;
        RECT  2.025 0.545 2.255 3.510 ;
        RECT  2.025 3.210 2.960 3.510 ;
        RECT  4.180 1.875 4.410 2.460 ;
        RECT  2.485 2.120 4.410 2.460 ;
        RECT  2.485 1.085 2.770 2.980 ;
        RECT  4.875 0.430 5.385 0.770 ;
        RECT  5.100 0.430 5.385 2.950 ;
        RECT  5.635 1.650 6.830 1.990 ;
        RECT  6.545 1.070 6.830 2.750 ;
        RECT  7.955 0.540 11.190 0.820 ;
        RECT  4.365 1.085 4.870 1.645 ;
        RECT  3.360 1.415 4.870 1.645 ;
        RECT  3.360 1.415 3.705 1.890 ;
        RECT  9.905 1.710 11.235 2.040 ;
        RECT  9.905 1.710 10.245 2.770 ;
        RECT  7.275 2.535 10.245 2.770 ;
        RECT  4.640 1.085 4.870 3.410 ;
        RECT  4.365 2.690 4.870 3.410 ;
        RECT  5.615 2.980 7.505 3.210 ;
        RECT  7.275 2.535 7.505 3.210 ;
        RECT  4.365 3.180 5.845 3.410 ;
        RECT  7.245 0.515 7.585 1.355 ;
        RECT  7.245 1.100 12.050 1.355 ;
        RECT  11.765 1.100 12.050 3.255 ;
        RECT  7.960 3.025 12.050 3.255 ;
    END
END TLATNTSCA_X12_18_SVT_WB

MACRO TLATNSR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNSR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.820 3.270 2.100 ;
        RECT  2.520 1.820 2.860 2.250 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.424  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.695 2.505 3.535 2.735 ;
        RECT  3.180 2.400 3.535 2.735 ;
        RECT  0.695 2.025 1.225 2.735 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.220 2.330 10.860 3.295 ;
        RECT  10.630 0.575 10.860 3.295 ;
        RECT  10.575 0.575 10.860 1.445 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.930 2.380 9.340 2.705 ;
        RECT  9.000 0.630 9.340 2.705 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.163  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.810 2.210 2.270 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.690 2.105 6.245 2.660 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  11.215 2.375 11.600 4.100 ;
        RECT  9.730 3.570 10.145 4.100 ;
        RECT  6.395 3.570 6.735 4.100 ;
        RECT  4.935 2.965 5.165 4.100 ;
        RECT  0.995 3.515 1.225 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  11.210 -0.180 11.615 1.470 ;
        RECT  9.815 -0.180 10.045 0.875 ;
        RECT  6.915 -0.180 7.225 1.430 ;
        RECT  5.105 -0.180 5.335 1.240 ;
        RECT  1.565 -0.180 1.795 1.035 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.550 0.775 1.015 1.580 ;
        RECT  0.235 1.340 1.015 1.580 ;
        RECT  0.235 1.350 4.135 1.580 ;
        RECT  3.905 1.350 4.135 2.730 ;
        RECT  0.235 1.340 0.465 3.430 ;
        RECT  3.445 0.705 4.595 1.045 ;
        RECT  4.365 2.335 5.440 2.675 ;
        RECT  4.365 0.705 4.595 3.305 ;
        RECT  1.665 2.965 4.595 3.305 ;
        RECT  4.825 1.645 6.685 1.875 ;
        RECT  6.255 0.980 6.685 1.875 ;
        RECT  4.825 1.645 5.055 2.005 ;
        RECT  6.475 1.780 7.210 2.120 ;
        RECT  6.475 1.780 6.705 3.285 ;
        RECT  5.690 2.945 6.705 3.285 ;
        RECT  7.470 1.100 7.940 1.440 ;
        RECT  9.670 1.740 10.400 2.085 ;
        RECT  7.470 1.100 7.700 3.285 ;
        RECT  7.210 2.845 7.700 3.285 ;
        RECT  9.670 1.740 9.900 3.285 ;
        RECT  7.210 3.035 9.900 3.285 ;
    END
END TLATNSR_X4_18_SVT_WB

MACRO TLATNSR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNSR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.820 3.270 2.100 ;
        RECT  2.520 1.820 2.860 2.250 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.291  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.695 2.505 3.530 2.735 ;
        RECT  3.185 2.400 3.530 2.735 ;
        RECT  0.695 2.280 1.000 2.735 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.610 2.365 10.195 3.295 ;
        RECT  9.965 0.575 10.195 3.295 ;
        RECT  9.910 0.575 10.195 1.445 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.930 2.380 8.675 2.705 ;
        RECT  8.335 0.630 8.675 2.705 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.810 2.210 2.270 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.690 2.105 6.245 2.660 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.065 3.570 9.480 4.100 ;
        RECT  6.395 3.570 6.735 4.100 ;
        RECT  4.935 2.965 5.165 4.100 ;
        RECT  0.995 3.515 1.225 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.150 -0.180 9.380 0.875 ;
        RECT  5.105 -0.180 5.335 1.240 ;
        RECT  1.565 -0.180 1.795 1.035 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.585 0.750 0.970 1.580 ;
        RECT  0.235 1.350 4.135 1.580 ;
        RECT  3.905 1.350 4.135 2.730 ;
        RECT  0.235 1.350 0.465 3.430 ;
        RECT  3.445 0.705 4.595 1.045 ;
        RECT  4.365 2.335 5.440 2.675 ;
        RECT  4.365 0.705 4.595 3.305 ;
        RECT  1.665 2.965 4.595 3.305 ;
        RECT  4.825 1.645 6.685 1.875 ;
        RECT  6.255 0.980 6.685 1.875 ;
        RECT  4.825 1.645 5.055 2.005 ;
        RECT  6.475 1.780 7.210 2.120 ;
        RECT  6.475 1.780 6.705 3.285 ;
        RECT  5.690 2.945 6.705 3.285 ;
        RECT  7.470 1.100 7.940 1.440 ;
        RECT  9.080 1.740 9.735 2.130 ;
        RECT  7.470 1.100 7.700 3.285 ;
        RECT  7.210 2.845 7.700 3.285 ;
        RECT  9.080 1.740 9.370 3.285 ;
        RECT  7.210 3.035 9.370 3.285 ;
    END
END TLATNSR_X2_18_SVT_WB

MACRO TLATNSR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNSR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.820 3.270 2.100 ;
        RECT  2.520 1.820 2.860 2.250 ;
        END
    END D
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.291  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.825 2.505 3.555 2.735 ;
        RECT  3.175 2.400 3.555 2.735 ;
        RECT  0.825 2.315 1.540 2.735 ;
        END
    END GN
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.610 2.365 10.195 2.665 ;
        RECT  9.965 0.575 10.195 2.665 ;
        RECT  9.910 0.575 10.195 0.915 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.930 2.380 8.675 2.705 ;
        RECT  8.335 0.630 8.675 2.705 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.132  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.810 2.210 2.270 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.169  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.690 2.105 6.245 2.660 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.065 3.570 9.480 4.100 ;
        RECT  6.395 3.570 6.735 4.100 ;
        RECT  4.935 2.965 5.165 4.100 ;
        RECT  0.995 3.515 1.225 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.150 -0.180 9.380 0.875 ;
        RECT  6.945 -0.180 7.240 1.495 ;
        RECT  5.105 -0.180 5.335 1.240 ;
        RECT  1.565 -0.180 1.795 1.035 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.595 0.775 0.985 1.580 ;
        RECT  0.235 1.325 0.985 1.580 ;
        RECT  0.235 1.350 4.135 1.580 ;
        RECT  3.905 1.350 4.135 2.730 ;
        RECT  0.235 1.325 0.465 3.430 ;
        RECT  3.445 0.705 4.595 1.045 ;
        RECT  4.365 2.335 5.440 2.675 ;
        RECT  4.365 0.705 4.595 3.305 ;
        RECT  1.665 2.965 4.595 3.305 ;
        RECT  4.825 1.645 6.685 1.875 ;
        RECT  6.255 0.980 6.685 1.875 ;
        RECT  4.825 1.645 5.055 2.005 ;
        RECT  6.475 1.780 7.210 2.120 ;
        RECT  6.475 1.780 6.705 3.285 ;
        RECT  5.690 2.945 6.705 3.285 ;
        RECT  7.470 1.100 7.940 1.440 ;
        RECT  9.080 1.105 9.735 1.495 ;
        RECT  7.470 1.100 7.700 3.285 ;
        RECT  7.210 2.845 7.700 3.285 ;
        RECT  9.080 1.105 9.370 3.285 ;
        RECT  7.210 3.035 9.370 3.285 ;
    END
END TLATNSR_X1_18_SVT_WB

MACRO TLATNCA_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.480  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.245 1.680 7.025 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.705 0.840 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.371  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.030 1.725 10.435 3.410 ;
        RECT  10.060 0.540 10.435 3.410 ;
        RECT  8.660 1.725 10.435 2.175 ;
        RECT  8.660 0.490 9.170 3.445 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  9.400 2.635 9.690 4.100 ;
        RECT  5.240 3.440 6.050 4.100 ;
        RECT  2.810 2.690 3.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  9.400 -0.180 9.690 1.300 ;
        RECT  4.990 -0.180 5.330 0.420 ;
        RECT  2.810 -0.180 3.150 1.375 ;
        RECT  0.235 -0.180 0.935 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.255 0.545 1.485 3.510 ;
        RECT  1.255 3.210 2.190 3.510 ;
        RECT  1.715 2.120 3.575 2.460 ;
        RECT  1.715 1.085 2.000 2.980 ;
        RECT  4.040 0.460 4.550 0.835 ;
        RECT  4.265 0.460 4.550 2.950 ;
        RECT  4.800 1.650 5.995 1.990 ;
        RECT  5.710 1.085 5.995 2.750 ;
        RECT  3.530 1.085 3.870 1.890 ;
        RECT  2.590 1.605 4.035 1.890 ;
        RECT  7.465 1.710 7.805 2.875 ;
        RECT  6.820 2.535 7.805 2.875 ;
        RECT  3.805 1.555 4.035 3.410 ;
        RECT  3.530 2.690 4.035 3.410 ;
        RECT  4.780 2.980 7.050 3.210 ;
        RECT  6.820 2.535 7.050 3.210 ;
        RECT  3.530 3.180 5.010 3.410 ;
        RECT  6.410 0.515 6.750 1.355 ;
        RECT  6.410 1.100 8.430 1.355 ;
        RECT  8.145 1.100 8.430 3.445 ;
        RECT  7.280 3.105 8.430 3.445 ;
    END
END TLATNCA_X8_18_SVT_WB

MACRO TLATNCA_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.480  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.225 1.680 6.960 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.705 0.840 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.239  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.120 2.480 10.465 3.445 ;
        RECT  8.660 1.125 10.465 1.360 ;
        RECT  10.120 0.490 10.465 1.360 ;
        RECT  8.660 2.480 10.465 2.740 ;
        RECT  9.495 1.125 9.940 2.740 ;
        RECT  8.660 2.480 9.040 3.460 ;
        RECT  8.660 0.490 9.035 1.360 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.430 3.045 9.740 4.100 ;
        RECT  5.240 3.440 6.050 4.100 ;
        RECT  2.810 2.690 3.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.390 -0.180 9.730 0.845 ;
        RECT  4.990 -0.180 5.330 0.425 ;
        RECT  2.810 -0.180 3.150 1.375 ;
        RECT  0.235 -0.180 0.935 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.255 0.545 1.485 3.510 ;
        RECT  1.255 3.210 2.190 3.510 ;
        RECT  1.715 2.120 3.575 2.460 ;
        RECT  1.715 1.085 2.000 2.980 ;
        RECT  4.040 0.490 4.550 0.845 ;
        RECT  4.265 0.490 4.550 2.950 ;
        RECT  4.800 1.650 5.995 1.990 ;
        RECT  5.710 1.085 5.995 2.750 ;
        RECT  3.530 1.085 3.870 1.890 ;
        RECT  2.590 1.605 4.035 1.890 ;
        RECT  7.465 1.770 7.805 2.875 ;
        RECT  6.820 2.535 7.805 2.875 ;
        RECT  3.805 1.555 4.035 3.410 ;
        RECT  3.530 2.690 4.035 3.410 ;
        RECT  4.780 2.980 7.050 3.210 ;
        RECT  6.820 2.535 7.050 3.210 ;
        RECT  3.530 3.180 5.010 3.410 ;
        RECT  6.410 0.565 6.765 1.380 ;
        RECT  6.410 1.110 8.430 1.380 ;
        RECT  8.180 1.670 8.965 1.910 ;
        RECT  8.180 1.110 8.430 3.445 ;
        RECT  7.280 3.105 8.430 3.445 ;
    END
END TLATNCA_X6_18_SVT_WB

MACRO TLATNCA_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.505 1.210 7.140 1.760 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.705 1.050 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.310 0.490 8.820 3.445 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  9.050 2.635 9.340 4.100 ;
        RECT  5.450 3.440 6.260 4.100 ;
        RECT  3.020 2.690 3.360 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  9.050 -0.180 9.340 1.300 ;
        RECT  5.200 -0.180 5.540 0.820 ;
        RECT  3.020 -0.180 3.360 1.375 ;
        RECT  0.445 -0.180 1.145 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.465 0.545 1.695 3.510 ;
        RECT  1.465 3.210 2.400 3.510 ;
        RECT  1.925 2.120 3.785 2.460 ;
        RECT  1.925 1.085 2.210 2.980 ;
        RECT  4.250 0.560 4.760 0.900 ;
        RECT  4.475 0.560 4.760 2.950 ;
        RECT  5.010 1.650 6.205 1.990 ;
        RECT  5.920 1.130 6.205 2.750 ;
        RECT  3.740 1.085 4.080 1.890 ;
        RECT  2.800 1.605 4.245 1.890 ;
        RECT  7.080 2.095 7.420 2.875 ;
        RECT  6.435 2.535 7.420 2.875 ;
        RECT  4.015 1.555 4.245 3.410 ;
        RECT  3.740 2.690 4.245 3.410 ;
        RECT  4.990 2.980 6.665 3.210 ;
        RECT  6.435 2.535 6.665 3.210 ;
        RECT  3.740 3.180 5.220 3.410 ;
        RECT  6.000 0.430 8.080 0.770 ;
        RECT  7.795 0.430 8.080 3.445 ;
        RECT  6.895 3.105 8.080 3.445 ;
    END
END TLATNCA_X4_18_SVT_WB

MACRO TLATNCA_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.730 1.660 6.020 2.360 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.540 0.540 2.265 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.899  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.335 0.815 7.700 2.980 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  4.790 3.445 5.545 4.100 ;
        RECT  2.340 2.525 2.680 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  6.600 -0.180 6.940 0.835 ;
        RECT  4.520 -0.180 4.860 0.820 ;
        RECT  2.340 -0.180 2.680 1.210 ;
        RECT  0.180 -0.180 0.520 0.485 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.770 0.410 1.290 0.690 ;
        RECT  0.770 0.410 1.000 3.370 ;
        RECT  0.770 3.045 1.770 3.370 ;
        RECT  1.230 1.955 3.070 2.295 ;
        RECT  1.230 0.920 1.530 2.815 ;
        RECT  3.570 0.425 4.065 0.765 ;
        RECT  3.760 0.425 4.065 1.460 ;
        RECT  3.760 0.425 3.990 3.050 ;
        RECT  3.760 2.735 4.100 3.050 ;
        RECT  5.135 1.135 5.495 1.635 ;
        RECT  4.220 1.635 5.365 1.995 ;
        RECT  5.080 1.635 5.365 2.755 ;
        RECT  3.060 0.920 3.400 1.725 ;
        RECT  2.120 1.440 3.530 1.725 ;
        RECT  5.595 2.590 6.500 2.880 ;
        RECT  5.595 2.590 5.825 3.215 ;
        RECT  4.330 2.985 5.825 3.215 ;
        RECT  3.300 1.440 3.530 3.510 ;
        RECT  3.060 2.525 3.530 3.510 ;
        RECT  4.330 2.985 4.560 3.510 ;
        RECT  3.060 3.280 4.560 3.510 ;
        RECT  5.220 0.435 5.955 0.775 ;
        RECT  5.725 0.435 5.955 1.430 ;
        RECT  5.725 1.200 7.105 1.430 ;
        RECT  6.820 1.200 7.105 3.450 ;
        RECT  6.055 3.110 7.105 3.450 ;
    END
END TLATNCA_X3_18_SVT_WB

MACRO TLATNCA_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.730 1.450 6.020 2.235 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.540 0.540 2.710 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.054  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.335 0.470 7.700 3.450 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  4.790 3.445 5.545 4.100 ;
        RECT  2.340 2.525 2.680 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  6.650 -0.180 6.940 0.810 ;
        RECT  4.520 -0.180 4.860 0.875 ;
        RECT  2.340 -0.180 2.680 1.210 ;
        RECT  0.180 -0.180 0.520 0.485 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.770 0.410 1.290 0.690 ;
        RECT  0.770 0.410 1.000 3.370 ;
        RECT  0.770 3.045 1.770 3.370 ;
        RECT  1.230 1.955 3.070 2.295 ;
        RECT  1.230 0.920 1.530 2.815 ;
        RECT  3.570 0.435 4.090 0.775 ;
        RECT  3.760 0.435 4.090 1.475 ;
        RECT  3.760 0.435 3.990 3.050 ;
        RECT  3.760 2.735 4.100 3.050 ;
        RECT  5.080 1.135 5.500 1.475 ;
        RECT  4.220 1.675 5.365 2.015 ;
        RECT  5.080 1.135 5.365 2.755 ;
        RECT  3.060 0.935 3.400 1.725 ;
        RECT  2.120 1.440 3.530 1.725 ;
        RECT  5.595 2.590 6.500 2.880 ;
        RECT  5.595 2.590 5.825 3.215 ;
        RECT  4.330 2.985 5.825 3.215 ;
        RECT  3.300 1.440 3.530 3.510 ;
        RECT  3.060 2.525 3.530 3.510 ;
        RECT  4.330 2.985 4.560 3.510 ;
        RECT  3.060 3.280 4.560 3.510 ;
        RECT  5.220 0.430 6.420 0.770 ;
        RECT  6.190 0.430 6.420 1.290 ;
        RECT  6.190 1.060 7.105 1.290 ;
        RECT  6.810 1.060 7.105 3.450 ;
        RECT  6.055 3.110 7.105 3.450 ;
    END
END TLATNCA_X2_18_SVT_WB

MACRO TLATNCA_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.310 1.680 8.525 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.705 0.840 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.926  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.000 0.490 17.340 3.355 ;
        RECT  11.510 1.725 17.340 2.170 ;
        RECT  15.680 0.555 16.020 3.355 ;
        RECT  14.240 0.570 14.580 3.410 ;
        RECT  12.880 1.725 13.285 3.410 ;
        RECT  12.910 0.540 13.285 3.410 ;
        RECT  11.510 1.725 13.285 2.175 ;
        RECT  11.510 1.725 11.890 3.445 ;
        RECT  11.510 0.490 11.880 3.445 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 18.480 4.100 ;
        RECT  17.720 2.565 18.060 4.100 ;
        RECT  14.960 2.495 15.300 4.100 ;
        RECT  12.200 2.635 12.540 4.100 ;
        RECT  5.305 3.440 6.645 4.100 ;
        RECT  2.810 2.690 3.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 18.480 0.180 ;
        RECT  17.720 -0.180 18.060 1.270 ;
        RECT  14.960 -0.180 15.300 1.285 ;
        RECT  12.200 -0.180 12.540 1.300 ;
        RECT  5.055 -0.180 5.395 0.415 ;
        RECT  2.875 -0.180 3.215 1.185 ;
        RECT  0.235 -0.180 0.935 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.255 0.545 1.485 3.510 ;
        RECT  1.255 3.210 2.190 3.510 ;
        RECT  3.410 1.875 3.640 2.460 ;
        RECT  1.715 2.120 3.640 2.460 ;
        RECT  1.715 1.085 2.000 2.980 ;
        RECT  4.105 0.430 4.615 0.770 ;
        RECT  4.330 0.430 4.615 2.950 ;
        RECT  4.865 1.650 6.060 1.990 ;
        RECT  5.775 1.070 6.060 2.750 ;
        RECT  7.185 0.540 10.420 0.820 ;
        RECT  3.595 1.085 4.100 1.645 ;
        RECT  2.590 1.415 4.100 1.645 ;
        RECT  2.590 1.415 2.935 1.890 ;
        RECT  9.135 1.710 10.465 2.040 ;
        RECT  9.135 1.710 9.475 2.770 ;
        RECT  6.505 2.535 9.475 2.770 ;
        RECT  3.870 1.085 4.100 3.410 ;
        RECT  3.595 2.690 4.100 3.410 ;
        RECT  4.845 2.980 6.735 3.210 ;
        RECT  6.505 2.535 6.735 3.210 ;
        RECT  3.595 3.180 5.075 3.410 ;
        RECT  6.475 0.515 6.815 1.355 ;
        RECT  6.475 1.100 11.280 1.355 ;
        RECT  10.995 1.100 11.280 3.255 ;
        RECT  7.190 3.025 11.280 3.255 ;
    END
END TLATNCA_X20_18_SVT_WB

MACRO TLATNCA_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.310 1.680 8.525 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.705 0.840 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.741  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.680 0.555 16.020 3.355 ;
        RECT  11.510 1.725 16.020 2.170 ;
        RECT  14.240 0.570 14.580 3.410 ;
        RECT  12.880 1.725 13.285 3.410 ;
        RECT  12.910 0.540 13.285 3.410 ;
        RECT  11.510 1.725 13.285 2.175 ;
        RECT  11.510 1.725 11.890 3.445 ;
        RECT  11.510 0.490 11.880 3.445 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.800 4.100 ;
        RECT  14.960 2.495 15.300 4.100 ;
        RECT  12.200 2.635 12.540 4.100 ;
        RECT  5.305 3.440 6.645 4.100 ;
        RECT  2.810 2.690 3.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.800 0.180 ;
        RECT  14.960 -0.180 15.300 1.285 ;
        RECT  12.200 -0.180 12.540 1.300 ;
        RECT  5.055 -0.180 5.395 0.415 ;
        RECT  2.875 -0.180 3.215 1.185 ;
        RECT  0.235 -0.180 0.935 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.255 0.545 1.485 3.510 ;
        RECT  1.255 3.210 2.190 3.510 ;
        RECT  3.410 1.875 3.640 2.460 ;
        RECT  1.715 2.120 3.640 2.460 ;
        RECT  1.715 1.085 2.000 2.980 ;
        RECT  4.105 0.430 4.615 0.770 ;
        RECT  4.330 0.430 4.615 2.950 ;
        RECT  4.865 1.650 6.060 1.990 ;
        RECT  5.775 1.070 6.060 2.750 ;
        RECT  7.185 0.540 10.420 0.820 ;
        RECT  3.595 1.085 4.100 1.645 ;
        RECT  2.590 1.415 4.100 1.645 ;
        RECT  2.590 1.415 2.935 1.890 ;
        RECT  9.135 1.710 10.465 2.040 ;
        RECT  9.135 1.710 9.475 2.770 ;
        RECT  6.505 2.535 9.475 2.770 ;
        RECT  3.870 1.085 4.100 3.410 ;
        RECT  3.595 2.690 4.100 3.410 ;
        RECT  4.845 2.980 6.735 3.210 ;
        RECT  6.505 2.535 6.735 3.210 ;
        RECT  3.595 3.180 5.075 3.410 ;
        RECT  6.475 0.515 6.815 1.355 ;
        RECT  6.475 1.100 11.280 1.355 ;
        RECT  10.995 1.100 11.280 3.255 ;
        RECT  7.190 3.025 11.280 3.255 ;
    END
END TLATNCA_X16_18_SVT_WB

MACRO TLATNCA_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN TLATNCA_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.270  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.310 1.680 8.525 2.230 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.705 0.840 2.660 ;
        END
    END E
    PIN ECK
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.556  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.360 0.570 14.700 3.410 ;
        RECT  11.510 1.725 14.700 2.170 ;
        RECT  12.880 1.725 13.285 3.410 ;
        RECT  12.910 0.540 13.285 3.410 ;
        RECT  11.510 1.725 13.285 2.175 ;
        RECT  11.510 1.725 11.890 3.445 ;
        RECT  11.510 0.490 11.880 3.445 ;
        END
    END ECK
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  15.080 2.495 15.420 4.100 ;
        RECT  13.640 2.600 13.980 4.100 ;
        RECT  12.200 2.635 12.540 4.100 ;
        RECT  5.305 3.440 6.645 4.100 ;
        RECT  2.810 2.690 3.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  15.080 -0.180 15.420 1.285 ;
        RECT  13.640 -0.180 13.980 1.295 ;
        RECT  12.200 -0.180 12.540 1.300 ;
        RECT  5.055 -0.180 5.395 0.415 ;
        RECT  2.875 -0.180 3.215 1.185 ;
        RECT  0.235 -0.180 0.935 0.515 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.255 0.545 1.485 3.510 ;
        RECT  1.255 3.210 2.190 3.510 ;
        RECT  3.410 1.875 3.640 2.460 ;
        RECT  1.715 2.120 3.640 2.460 ;
        RECT  1.715 1.085 2.000 2.980 ;
        RECT  4.105 0.430 4.615 0.770 ;
        RECT  4.330 0.430 4.615 2.950 ;
        RECT  4.865 1.650 6.060 1.990 ;
        RECT  5.775 1.070 6.060 2.750 ;
        RECT  7.185 0.540 10.420 0.820 ;
        RECT  3.595 1.085 4.100 1.645 ;
        RECT  2.590 1.415 4.100 1.645 ;
        RECT  2.590 1.415 2.935 1.890 ;
        RECT  9.135 1.710 10.465 2.040 ;
        RECT  9.135 1.710 9.475 2.770 ;
        RECT  6.505 2.535 9.475 2.770 ;
        RECT  3.870 1.085 4.100 3.410 ;
        RECT  3.595 2.690 4.100 3.410 ;
        RECT  4.845 2.980 6.735 3.210 ;
        RECT  6.505 2.535 6.735 3.210 ;
        RECT  3.595 3.180 5.075 3.410 ;
        RECT  6.475 0.515 6.815 1.355 ;
        RECT  6.475 1.100 11.280 1.355 ;
        RECT  10.995 1.100 11.280 3.255 ;
        RECT  7.190 3.025 11.280 3.255 ;
    END
END TLATNCA_X12_18_SVT_WB

MACRO TIEL_18_SVT_WB
    CLASS CORE ;
    FOREIGN TIEL_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.252  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.210 0.780 1.590 ;
        RECT  0.440 0.920 0.780 1.590 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  1.160 2.680 1.500 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  1.160 -0.180 1.500 1.235 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.440 2.160 0.780 3.070 ;
    END
END TIEL_18_SVT_WB

MACRO TIEH_18_SVT_WB
    CLASS CORE ;
    FOREIGN TIEH_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.276  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.440 2.815 0.980 3.270 ;
        RECT  0.440 2.605 0.750 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  1.210 2.815 1.500 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  1.160 -0.180 1.500 1.180 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.460 0.840 0.800 1.700 ;
    END
END TIEH_18_SVT_WB

MACRO SDFF_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFF_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.480 0.600 13.860 3.480 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.715 2.420 11.385 2.760 ;
        RECT  11.105 1.135 11.385 2.760 ;
        RECT  10.660 1.135 11.385 1.540 ;
        RECT  10.715 2.420 11.100 3.420 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.560 4.100 ;
        RECT  12.705 3.515 13.075 4.100 ;
        RECT  9.790 3.485 10.245 4.100 ;
        RECT  7.215 2.695 7.555 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.560 0.180 ;
        RECT  12.705 -0.180 13.060 0.405 ;
        RECT  9.900 -0.180 10.250 0.405 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.550 1.040 1.915 1.345 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.430 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  5.350 0.880 5.730 1.230 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.380 0.880 5.730 3.335 ;
        RECT  2.375 3.105 5.730 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.650 1.220 ;
        RECT  7.390 0.880 7.650 1.740 ;
        RECT  7.390 1.400 7.730 1.740 ;
        RECT  6.385 0.880 6.615 2.995 ;
        RECT  6.065 2.655 6.615 2.995 ;
        RECT  7.880 0.880 8.260 1.220 ;
        RECT  6.975 2.125 8.260 2.465 ;
        RECT  7.960 0.880 8.260 3.020 ;
        RECT  7.935 2.125 8.260 3.020 ;
        RECT  4.890 0.410 9.335 0.650 ;
        RECT  4.890 0.410 5.120 1.345 ;
        RECT  4.470 1.055 5.120 1.345 ;
        RECT  4.470 1.870 4.895 2.245 ;
        RECT  9.105 0.410 9.335 2.500 ;
        RECT  8.950 2.160 9.335 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  8.490 0.880 8.875 1.220 ;
        RECT  10.255 1.865 10.760 2.190 ;
        RECT  8.490 0.880 8.720 3.020 ;
        RECT  10.255 1.865 10.485 3.020 ;
        RECT  8.490 2.730 10.485 3.020 ;
        RECT  11.920 0.430 12.260 0.905 ;
        RECT  9.565 0.635 13.200 0.905 ;
        RECT  9.565 0.635 9.945 2.065 ;
        RECT  12.935 0.635 13.200 3.285 ;
        RECT  11.945 3.055 13.200 3.285 ;
        RECT  11.945 3.055 12.285 3.465 ;
    END
END SDFF_X4_18_SVT_WB

MACRO SDFF_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFF_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.920 0.600 13.300 3.480 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.990 1.135 11.220 2.760 ;
        RECT  10.715 2.420 11.100 3.420 ;
        RECT  10.660 1.135 11.220 1.540 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 13.440 4.100 ;
        RECT  12.145 3.515 12.515 4.100 ;
        RECT  9.790 3.485 10.245 4.100 ;
        RECT  7.215 2.695 7.555 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 13.440 0.180 ;
        RECT  12.145 -0.180 12.500 0.405 ;
        RECT  9.900 -0.180 10.250 0.405 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.550 1.040 1.915 1.345 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.430 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  5.350 0.880 5.730 1.230 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.380 0.880 5.730 3.335 ;
        RECT  2.375 3.105 5.730 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.650 1.220 ;
        RECT  7.390 0.880 7.650 1.740 ;
        RECT  7.390 1.400 7.730 1.740 ;
        RECT  6.385 0.880 6.615 2.995 ;
        RECT  6.065 2.655 6.615 2.995 ;
        RECT  7.880 0.880 8.260 1.220 ;
        RECT  6.975 2.125 8.260 2.465 ;
        RECT  7.960 0.880 8.260 3.020 ;
        RECT  7.935 2.125 8.260 3.020 ;
        RECT  4.890 0.410 9.335 0.650 ;
        RECT  4.890 0.410 5.120 1.345 ;
        RECT  4.470 1.055 5.120 1.345 ;
        RECT  4.470 1.870 4.895 2.245 ;
        RECT  9.105 0.410 9.335 2.500 ;
        RECT  8.950 2.160 9.335 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  8.490 0.880 8.875 1.220 ;
        RECT  10.255 1.865 10.760 2.190 ;
        RECT  8.490 0.880 8.720 3.020 ;
        RECT  10.255 1.865 10.485 3.020 ;
        RECT  8.490 2.730 10.485 3.020 ;
        RECT  11.360 0.430 11.700 0.905 ;
        RECT  9.565 0.635 12.640 0.905 ;
        RECT  9.565 0.635 9.945 2.065 ;
        RECT  12.375 0.635 12.640 3.285 ;
        RECT  11.385 3.055 12.640 3.285 ;
        RECT  11.385 3.055 11.725 3.465 ;
    END
END SDFF_X2_18_SVT_WB

MACRO SDFF_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFF_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.920 0.515 13.300 3.480 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.990 1.135 11.220 2.760 ;
        RECT  10.715 2.420 11.100 3.370 ;
        RECT  10.660 1.135 11.220 1.540 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 13.440 4.100 ;
        RECT  12.145 3.515 12.515 4.100 ;
        RECT  9.790 3.485 10.245 4.100 ;
        RECT  7.215 2.695 7.555 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 13.440 0.180 ;
        RECT  12.145 -0.180 12.500 0.405 ;
        RECT  9.900 -0.180 10.250 0.405 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.550 1.040 1.915 1.345 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.430 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  5.350 0.880 5.730 1.230 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.380 0.880 5.730 3.335 ;
        RECT  2.375 3.105 5.730 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.650 1.220 ;
        RECT  7.390 0.880 7.650 1.740 ;
        RECT  7.390 1.400 7.730 1.740 ;
        RECT  6.385 0.880 6.615 2.995 ;
        RECT  6.065 2.655 6.615 2.995 ;
        RECT  7.880 0.880 8.260 1.220 ;
        RECT  6.975 2.125 8.260 2.465 ;
        RECT  7.960 0.880 8.260 3.020 ;
        RECT  7.935 2.125 8.260 3.020 ;
        RECT  4.890 0.410 9.335 0.650 ;
        RECT  4.890 0.410 5.120 1.345 ;
        RECT  4.470 1.055 5.120 1.345 ;
        RECT  4.470 1.870 4.895 2.245 ;
        RECT  9.105 0.410 9.335 2.500 ;
        RECT  8.950 2.160 9.335 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  8.490 0.880 8.875 1.220 ;
        RECT  10.255 1.865 10.760 2.190 ;
        RECT  8.490 0.880 8.720 3.020 ;
        RECT  10.255 1.865 10.485 3.020 ;
        RECT  8.490 2.730 10.485 3.020 ;
        RECT  11.360 0.430 11.700 0.905 ;
        RECT  9.565 0.635 12.640 0.905 ;
        RECT  9.565 0.635 9.945 2.065 ;
        RECT  12.375 0.635 12.640 3.285 ;
        RECT  11.385 3.055 12.640 3.285 ;
        RECT  11.385 3.055 11.725 3.465 ;
    END
END SDFF_X1_18_SVT_WB

MACRO SDFFTR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFTR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.305 1.595 6.085 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.311  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 1.705 5.005 2.270 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.625 0.470 16.120 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.800 2.480 13.445 2.775 ;
        RECT  13.215 1.145 13.445 2.775 ;
        RECT  12.800 1.145 13.445 1.570 ;
        RECT  12.800 2.480 13.180 3.255 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.095 3.460 1.590 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.915 2.185 2.150 ;
        RECT  1.900 1.765 2.185 2.150 ;
        RECT  0.125 1.915 1.000 2.255 ;
        RECT  0.125 1.655 0.430 2.255 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.665 1.210 1.440 1.590 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.800 4.100 ;
        RECT  15.000 3.110 15.340 4.100 ;
        RECT  12.065 3.485 12.405 4.100 ;
        RECT  9.665 2.700 10.005 4.100 ;
        RECT  5.910 3.370 6.250 4.100 ;
        RECT  4.050 3.560 4.390 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.800 0.180 ;
        RECT  15.000 -0.180 15.340 0.810 ;
        RECT  12.180 -0.180 12.520 0.455 ;
        RECT  5.980 -0.180 6.320 0.360 ;
        RECT  4.810 -0.180 5.150 0.355 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.575 0.520 0.915 ;
        RECT  0.180 0.635 1.900 0.915 ;
        RECT  1.670 0.635 1.900 1.435 ;
        RECT  1.670 1.095 2.655 1.435 ;
        RECT  1.910 2.435 2.655 2.720 ;
        RECT  2.415 1.095 2.655 2.720 ;
        RECT  0.180 2.485 2.655 2.720 ;
        RECT  0.180 2.485 0.520 3.295 ;
        RECT  3.345 2.930 3.755 3.320 ;
        RECT  3.345 3.090 5.195 3.320 ;
        RECT  4.795 3.090 5.195 3.460 ;
        RECT  5.350 1.090 6.545 1.365 ;
        RECT  6.315 1.090 6.545 2.750 ;
        RECT  5.350 2.465 6.545 2.750 ;
        RECT  2.130 0.520 2.470 0.860 ;
        RECT  2.130 0.620 7.725 0.850 ;
        RECT  2.130 0.620 3.990 0.860 ;
        RECT  3.760 0.620 3.990 2.400 ;
        RECT  2.885 2.170 3.990 2.400 ;
        RECT  7.480 0.620 7.725 2.720 ;
        RECT  2.885 2.170 3.115 3.280 ;
        RECT  2.065 3.005 3.115 3.280 ;
        RECT  8.415 1.450 10.190 1.790 ;
        RECT  8.415 0.930 8.730 2.720 ;
        RECT  10.190 0.930 10.670 1.220 ;
        RECT  9.420 2.130 10.670 2.470 ;
        RECT  10.420 0.930 10.670 3.020 ;
        RECT  10.385 2.130 10.670 3.020 ;
        RECT  7.955 0.410 11.685 0.700 ;
        RECT  11.425 0.410 11.685 2.500 ;
        RECT  7.955 0.410 8.185 3.390 ;
        RECT  6.775 1.080 7.080 3.390 ;
        RECT  7.955 2.880 8.220 3.390 ;
        RECT  6.775 3.160 8.220 3.390 ;
        RECT  12.700 1.800 12.985 2.250 ;
        RECT  11.915 2.020 12.985 2.250 ;
        RECT  10.910 0.930 11.195 3.020 ;
        RECT  11.915 2.020 12.145 3.020 ;
        RECT  10.910 2.730 12.145 3.020 ;
        RECT  14.200 0.470 14.555 0.915 ;
        RECT  12.140 0.685 14.555 0.915 ;
        RECT  12.140 0.685 12.370 1.790 ;
        RECT  11.915 1.450 12.370 1.790 ;
        RECT  14.325 1.860 15.395 2.200 ;
        RECT  14.325 0.470 14.555 3.450 ;
        RECT  14.200 3.110 14.555 3.450 ;
    END
END SDFFTR_X4_18_SVT_WB

MACRO SDFFTR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFTR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.305 1.595 6.085 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.311  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 1.705 5.005 2.270 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.065 0.470 15.540 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.215 1.145 13.445 2.775 ;
        RECT  12.905 2.480 13.320 3.340 ;
        RECT  12.800 1.145 13.445 1.570 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.095 3.460 1.590 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.915 2.185 2.150 ;
        RECT  1.900 1.765 2.185 2.150 ;
        RECT  0.125 1.915 1.000 2.255 ;
        RECT  0.125 1.655 0.430 2.255 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.665 1.210 1.440 1.590 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  14.440 3.110 14.780 4.100 ;
        RECT  12.065 3.485 12.405 4.100 ;
        RECT  9.665 2.700 10.005 4.100 ;
        RECT  5.910 3.370 6.250 4.100 ;
        RECT  4.050 3.560 4.390 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  14.440 -0.180 14.780 0.810 ;
        RECT  12.180 -0.180 12.520 0.455 ;
        RECT  5.980 -0.180 6.320 0.360 ;
        RECT  4.810 -0.180 5.150 0.355 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.575 0.520 0.915 ;
        RECT  0.180 0.635 1.900 0.915 ;
        RECT  1.670 0.635 1.900 1.435 ;
        RECT  1.670 1.095 2.655 1.435 ;
        RECT  1.910 2.435 2.655 2.720 ;
        RECT  2.415 1.095 2.655 2.720 ;
        RECT  0.180 2.485 2.655 2.720 ;
        RECT  0.180 2.485 0.520 3.295 ;
        RECT  3.345 2.930 3.755 3.320 ;
        RECT  3.345 3.090 5.195 3.320 ;
        RECT  4.795 3.090 5.195 3.460 ;
        RECT  5.350 1.090 6.545 1.365 ;
        RECT  6.315 1.090 6.545 2.750 ;
        RECT  5.350 2.465 6.545 2.750 ;
        RECT  2.130 0.520 2.470 0.860 ;
        RECT  2.130 0.620 7.725 0.850 ;
        RECT  2.130 0.620 3.990 0.860 ;
        RECT  3.760 0.620 3.990 2.400 ;
        RECT  2.885 2.170 3.990 2.400 ;
        RECT  7.480 0.620 7.725 2.720 ;
        RECT  2.885 2.170 3.115 3.280 ;
        RECT  2.065 3.005 3.115 3.280 ;
        RECT  8.415 1.450 10.190 1.790 ;
        RECT  8.415 0.930 8.730 2.720 ;
        RECT  10.190 0.930 10.670 1.220 ;
        RECT  9.420 2.130 10.670 2.470 ;
        RECT  10.420 0.930 10.670 3.020 ;
        RECT  10.385 2.130 10.670 3.020 ;
        RECT  7.955 0.410 11.685 0.700 ;
        RECT  11.425 0.410 11.685 2.500 ;
        RECT  7.955 0.410 8.185 3.390 ;
        RECT  6.775 1.080 7.080 3.390 ;
        RECT  7.955 2.880 8.220 3.390 ;
        RECT  6.775 3.160 8.220 3.390 ;
        RECT  12.700 1.800 12.985 2.250 ;
        RECT  11.915 2.020 12.985 2.250 ;
        RECT  10.910 0.930 11.195 3.020 ;
        RECT  11.915 2.020 12.145 3.020 ;
        RECT  10.910 2.730 12.145 3.020 ;
        RECT  13.640 0.470 13.995 0.915 ;
        RECT  12.140 0.685 13.995 0.915 ;
        RECT  12.140 0.685 12.370 1.790 ;
        RECT  11.915 1.450 12.370 1.790 ;
        RECT  13.765 1.860 14.835 2.200 ;
        RECT  13.765 0.470 13.995 3.450 ;
        RECT  13.640 3.110 13.995 3.450 ;
    END
END SDFFTR_X2_18_SVT_WB

MACRO SDFFTR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFTR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.305 1.595 6.085 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.311  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.230 1.705 5.005 2.270 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.065 0.470 15.540 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.215 1.145 13.445 2.775 ;
        RECT  12.905 2.480 13.320 3.340 ;
        RECT  12.800 1.145 13.445 1.570 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.905 1.095 3.460 1.590 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.915 2.185 2.150 ;
        RECT  1.900 1.765 2.185 2.150 ;
        RECT  0.125 1.915 1.000 2.255 ;
        RECT  0.125 1.655 0.430 2.255 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.665 1.210 1.440 1.590 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  14.440 3.110 14.780 4.100 ;
        RECT  12.065 3.485 12.405 4.100 ;
        RECT  9.665 2.700 10.005 4.100 ;
        RECT  5.910 3.370 6.250 4.100 ;
        RECT  4.050 3.560 4.390 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  14.440 -0.180 14.780 0.810 ;
        RECT  12.180 -0.180 12.520 0.455 ;
        RECT  5.980 -0.180 6.320 0.360 ;
        RECT  4.810 -0.180 5.150 0.355 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.575 0.520 0.915 ;
        RECT  0.180 0.635 1.900 0.915 ;
        RECT  1.670 0.635 1.900 1.435 ;
        RECT  1.670 1.095 2.655 1.435 ;
        RECT  1.910 2.435 2.655 2.720 ;
        RECT  2.415 1.095 2.655 2.720 ;
        RECT  0.180 2.485 2.655 2.720 ;
        RECT  0.180 2.485 0.520 3.295 ;
        RECT  3.345 2.930 3.755 3.320 ;
        RECT  3.345 3.090 5.195 3.320 ;
        RECT  4.795 3.090 5.195 3.460 ;
        RECT  5.350 1.090 6.545 1.365 ;
        RECT  6.315 1.090 6.545 2.750 ;
        RECT  5.350 2.465 6.545 2.750 ;
        RECT  2.130 0.520 2.470 0.860 ;
        RECT  2.130 0.620 7.725 0.850 ;
        RECT  2.130 0.620 3.990 0.860 ;
        RECT  3.760 0.620 3.990 2.400 ;
        RECT  2.885 2.170 3.990 2.400 ;
        RECT  7.480 0.620 7.725 2.720 ;
        RECT  2.885 2.170 3.115 3.280 ;
        RECT  2.065 3.005 3.115 3.280 ;
        RECT  8.415 1.450 10.190 1.790 ;
        RECT  8.415 0.930 8.730 2.720 ;
        RECT  10.190 0.930 10.670 1.220 ;
        RECT  9.420 2.130 10.670 2.470 ;
        RECT  10.420 0.930 10.670 3.020 ;
        RECT  10.385 2.130 10.670 3.020 ;
        RECT  7.955 0.410 11.685 0.700 ;
        RECT  11.425 0.410 11.685 2.500 ;
        RECT  7.955 0.410 8.185 3.390 ;
        RECT  6.775 1.080 7.080 3.390 ;
        RECT  7.955 2.880 8.220 3.390 ;
        RECT  6.775 3.160 8.220 3.390 ;
        RECT  12.700 1.800 12.985 2.250 ;
        RECT  11.915 2.020 12.985 2.250 ;
        RECT  10.910 0.930 11.195 3.020 ;
        RECT  11.915 2.020 12.145 3.020 ;
        RECT  10.910 2.730 12.145 3.020 ;
        RECT  13.640 0.470 13.995 0.915 ;
        RECT  12.140 0.685 13.995 0.915 ;
        RECT  12.140 0.685 12.370 1.790 ;
        RECT  11.915 1.450 12.370 1.790 ;
        RECT  13.765 1.860 14.835 2.200 ;
        RECT  13.765 0.470 13.995 3.450 ;
        RECT  13.640 3.110 13.995 3.450 ;
    END
END SDFFTR_X1_18_SVT_WB

MACRO SDFFS_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFS_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.035 1.045 15.555 3.410 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.505 2.505 17.220 2.815 ;
        RECT  16.920 1.045 17.220 2.815 ;
        RECT  16.505 1.045 17.220 1.400 ;
        RECT  16.505 2.505 16.830 3.405 ;
        RECT  16.505 0.575 16.830 1.400 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.805 1.750 12.195 2.305 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  17.210 3.050 17.550 4.100 ;
        RECT  15.820 2.575 16.110 4.100 ;
        RECT  14.285 3.430 14.635 4.100 ;
        RECT  11.890 3.570 13.170 4.100 ;
        RECT  7.750 3.530 9.030 4.100 ;
        RECT  3.855 3.570 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  17.210 -0.180 17.550 0.815 ;
        RECT  14.290 -0.180 14.630 0.350 ;
        RECT  12.460 -0.180 12.800 0.350 ;
        RECT  7.600 -0.180 7.940 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.535 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  5.770 0.940 6.120 1.310 ;
        RECT  5.870 0.940 6.120 2.995 ;
        RECT  4.985 2.705 6.120 2.995 ;
        RECT  4.010 1.055 4.240 3.340 ;
        RECT  2.375 3.105 4.240 3.340 ;
        RECT  4.985 2.705 5.215 3.340 ;
        RECT  2.375 3.110 5.215 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.500 1.045 7.080 1.385 ;
        RECT  6.850 2.090 8.460 2.350 ;
        RECT  6.850 1.045 7.080 2.840 ;
        RECT  6.500 2.555 7.080 2.840 ;
        RECT  7.450 1.565 9.075 1.860 ;
        RECT  8.790 1.045 9.075 2.840 ;
        RECT  8.735 1.565 9.075 2.840 ;
        RECT  8.735 2.500 9.910 2.840 ;
        RECT  8.310 2.580 9.910 2.840 ;
        RECT  6.660 3.070 10.080 3.300 ;
        RECT  5.455 3.270 7.100 3.510 ;
        RECT  9.795 3.070 10.080 3.510 ;
        RECT  5.100 0.410 7.100 0.640 ;
        RECT  6.725 0.585 11.110 0.815 ;
        RECT  5.100 0.410 5.330 1.350 ;
        RECT  4.470 1.120 5.330 1.350 ;
        RECT  9.305 0.585 9.535 1.905 ;
        RECT  9.305 1.565 9.620 1.905 ;
        RECT  10.770 0.585 11.110 2.305 ;
        RECT  4.470 2.015 5.525 2.395 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.765 1.045 10.155 1.385 ;
        RECT  10.030 1.180 10.540 1.615 ;
        RECT  13.185 2.005 13.565 2.365 ;
        RECT  10.310 1.180 10.540 3.340 ;
        RECT  10.310 2.530 10.630 3.340 ;
        RECT  13.185 2.005 13.415 3.340 ;
        RECT  10.310 3.105 13.415 3.340 ;
        RECT  12.505 1.045 14.585 1.360 ;
        RECT  12.505 1.045 12.765 1.995 ;
        RECT  14.250 1.045 14.585 2.945 ;
        RECT  13.645 2.595 14.585 2.945 ;
        RECT  13.645 2.595 13.910 3.425 ;
        RECT  11.600 0.585 16.275 0.815 ;
        RECT  11.600 0.585 11.860 1.385 ;
        RECT  11.345 1.025 11.860 1.385 ;
        RECT  16.040 0.585 16.275 1.960 ;
        RECT  11.345 1.025 11.575 2.875 ;
        RECT  11.010 2.535 12.610 2.875 ;
    END
END SDFFS_X4_18_SVT_WB

MACRO SDFFS_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFS_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.695 1.045 15.040 2.780 ;
        RECT  14.265 3.075 14.755 3.410 ;
        RECT  14.465 2.495 14.755 3.410 ;
        RECT  14.185 1.045 15.040 1.390 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.735 0.575 16.100 3.405 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.795 1.750 12.185 2.305 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  15.050 3.055 15.340 4.100 ;
        RECT  11.880 3.570 13.160 4.100 ;
        RECT  7.555 3.530 8.835 4.100 ;
        RECT  3.855 3.570 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  14.950 -0.180 15.320 0.350 ;
        RECT  12.450 -0.180 12.790 0.350 ;
        RECT  7.405 -0.180 7.745 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.535 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  5.575 0.940 5.925 1.310 ;
        RECT  5.675 0.940 5.925 2.995 ;
        RECT  4.930 2.705 5.925 2.995 ;
        RECT  4.010 1.055 4.240 3.340 ;
        RECT  2.375 3.105 4.240 3.340 ;
        RECT  4.930 2.705 5.160 3.340 ;
        RECT  2.375 3.110 5.160 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.305 1.045 6.885 1.385 ;
        RECT  6.655 2.090 8.265 2.350 ;
        RECT  6.655 1.045 6.885 2.840 ;
        RECT  6.305 2.555 6.885 2.840 ;
        RECT  7.255 1.565 8.880 1.860 ;
        RECT  8.595 1.045 8.880 2.840 ;
        RECT  8.540 1.565 8.880 2.840 ;
        RECT  8.540 2.500 9.715 2.840 ;
        RECT  8.115 2.580 9.715 2.840 ;
        RECT  6.465 3.070 9.885 3.300 ;
        RECT  5.390 3.270 6.905 3.510 ;
        RECT  9.600 3.070 9.885 3.510 ;
        RECT  5.100 0.410 6.905 0.640 ;
        RECT  6.530 0.585 10.915 0.815 ;
        RECT  5.100 0.410 5.330 1.350 ;
        RECT  4.470 1.120 5.330 1.350 ;
        RECT  9.110 0.585 9.340 1.905 ;
        RECT  9.110 1.565 9.425 1.905 ;
        RECT  4.470 1.055 4.755 2.295 ;
        RECT  4.470 1.915 5.320 2.295 ;
        RECT  10.575 0.585 10.915 2.305 ;
        RECT  4.470 1.055 4.700 2.875 ;
        RECT  9.570 1.045 9.960 1.385 ;
        RECT  9.835 1.180 10.345 1.615 ;
        RECT  13.175 2.005 13.490 2.365 ;
        RECT  10.115 1.180 10.345 3.340 ;
        RECT  10.115 2.530 10.435 3.340 ;
        RECT  13.175 2.005 13.405 3.340 ;
        RECT  10.115 3.105 13.405 3.340 ;
        RECT  12.495 1.045 13.950 1.360 ;
        RECT  12.495 1.045 12.755 1.995 ;
        RECT  13.720 1.645 14.235 1.995 ;
        RECT  13.720 1.045 13.950 3.425 ;
        RECT  13.635 2.595 13.950 3.425 ;
        RECT  11.590 0.585 15.505 0.815 ;
        RECT  11.590 0.585 11.850 1.385 ;
        RECT  11.220 1.025 11.850 1.385 ;
        RECT  15.270 0.585 15.505 1.960 ;
        RECT  11.220 1.025 11.565 2.875 ;
        RECT  10.815 2.535 12.600 2.875 ;
    END
END SDFFS_X2_18_SVT_WB

MACRO SDFFS_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFS_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.670 1.045 15.040 2.715 ;
        RECT  14.265 3.075 14.785 3.410 ;
        RECT  14.465 2.450 14.785 3.410 ;
        RECT  14.250 1.045 15.040 1.390 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.735 1.045 16.100 3.405 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.795 1.750 12.185 2.305 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  15.050 3.040 15.340 4.100 ;
        RECT  11.880 3.570 13.160 4.100 ;
        RECT  7.555 3.530 8.835 4.100 ;
        RECT  3.855 3.570 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  14.950 -0.180 15.320 0.350 ;
        RECT  12.450 -0.180 12.790 0.350 ;
        RECT  7.405 -0.180 7.745 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.535 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  5.575 0.940 5.925 1.310 ;
        RECT  5.675 0.940 5.925 2.995 ;
        RECT  4.930 2.705 5.925 2.995 ;
        RECT  4.010 1.055 4.240 3.340 ;
        RECT  2.375 3.105 4.240 3.340 ;
        RECT  4.930 2.705 5.160 3.340 ;
        RECT  2.375 3.110 5.160 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.305 1.045 6.885 1.385 ;
        RECT  6.655 2.090 8.265 2.350 ;
        RECT  6.655 1.045 6.885 2.840 ;
        RECT  6.305 2.555 6.885 2.840 ;
        RECT  7.255 1.565 8.880 1.860 ;
        RECT  8.595 1.045 8.880 2.840 ;
        RECT  8.540 1.565 8.880 2.840 ;
        RECT  8.540 2.500 9.715 2.840 ;
        RECT  8.115 2.580 9.715 2.840 ;
        RECT  6.465 3.070 9.885 3.300 ;
        RECT  5.390 3.270 6.905 3.510 ;
        RECT  9.600 3.070 9.885 3.510 ;
        RECT  5.100 0.410 6.905 0.640 ;
        RECT  6.530 0.585 10.915 0.815 ;
        RECT  5.100 0.410 5.330 1.350 ;
        RECT  4.470 1.055 5.330 1.350 ;
        RECT  9.110 0.585 9.340 1.905 ;
        RECT  9.110 1.565 9.425 1.905 ;
        RECT  4.470 1.055 4.755 2.365 ;
        RECT  10.575 0.585 10.915 2.305 ;
        RECT  4.470 1.985 5.285 2.365 ;
        RECT  4.470 1.055 4.700 2.875 ;
        RECT  9.570 1.045 9.960 1.385 ;
        RECT  9.835 1.180 10.345 1.615 ;
        RECT  13.175 2.005 13.555 2.300 ;
        RECT  10.115 1.180 10.345 3.340 ;
        RECT  10.115 2.530 10.435 3.340 ;
        RECT  13.175 2.005 13.405 3.340 ;
        RECT  10.115 3.105 13.405 3.340 ;
        RECT  12.495 1.045 14.015 1.360 ;
        RECT  12.495 1.045 12.755 1.995 ;
        RECT  13.785 1.645 14.235 1.995 ;
        RECT  13.785 1.045 14.015 2.875 ;
        RECT  13.635 2.530 14.015 2.875 ;
        RECT  11.590 0.585 15.505 0.815 ;
        RECT  11.590 0.585 11.850 1.385 ;
        RECT  11.240 1.025 11.850 1.385 ;
        RECT  15.270 0.585 15.505 1.960 ;
        RECT  11.240 1.025 11.565 2.875 ;
        RECT  10.815 2.535 12.600 2.875 ;
    END
END SDFFS_X1_18_SVT_WB

MACRO SDFFSR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFSR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.224  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.080 2.380 17.420 3.415 ;
        RECT  16.880 0.870 17.165 3.135 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.520 2.385 18.900 3.195 ;
        RECT  18.610 0.580 18.900 3.195 ;
        RECT  18.520 0.580 18.900 1.390 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.660 1.670 15.000 2.340 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.269  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.020 1.700 13.490 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 19.600 4.100 ;
        RECT  17.800 2.385 18.140 4.100 ;
        RECT  15.860 3.545 16.200 4.100 ;
        RECT  13.020 3.545 14.300 4.100 ;
        RECT  9.820 3.545 10.160 4.100 ;
        RECT  7.800 3.545 8.140 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 19.600 0.180 ;
        RECT  17.855 -0.180 18.140 1.390 ;
        RECT  14.140 -0.180 14.480 0.850 ;
        RECT  7.940 -0.180 8.280 0.815 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.610 1.100 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  4.430 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.635 1.725 0.870 ;
        RECT  0.470 0.635 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.455 0.970 5.685 3.335 ;
        RECT  2.375 3.105 5.685 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  7.040 2.565 8.700 2.855 ;
        RECT  6.375 0.970 6.715 1.310 ;
        RECT  6.485 1.505 9.100 1.765 ;
        RECT  8.760 1.505 9.100 1.845 ;
        RECT  6.485 0.970 6.715 2.855 ;
        RECT  6.375 2.515 6.715 2.855 ;
        RECT  7.230 1.995 7.570 2.335 ;
        RECT  7.230 2.105 10.220 2.335 ;
        RECT  9.935 0.970 10.220 2.855 ;
        RECT  9.060 2.105 10.220 2.855 ;
        RECT  9.060 2.515 10.865 2.855 ;
        RECT  11.095 1.960 11.410 2.300 ;
        RECT  11.095 1.960 11.325 3.315 ;
        RECT  6.560 3.085 11.325 3.315 ;
        RECT  6.560 3.085 6.900 3.425 ;
        RECT  4.890 0.410 7.285 0.640 ;
        RECT  9.365 0.410 12.330 0.740 ;
        RECT  6.945 0.410 7.285 1.275 ;
        RECT  9.365 0.410 9.705 1.275 ;
        RECT  6.945 1.045 9.705 1.275 ;
        RECT  4.890 0.410 5.120 1.335 ;
        RECT  4.470 1.055 5.120 1.335 ;
        RECT  10.450 0.410 10.705 1.830 ;
        RECT  12.100 0.410 12.330 2.100 ;
        RECT  4.470 1.840 5.095 2.235 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  10.935 0.970 11.225 1.310 ;
        RECT  10.935 1.035 11.870 1.310 ;
        RECT  11.640 1.035 11.870 3.315 ;
        RECT  11.555 2.515 11.870 3.315 ;
        RECT  15.690 2.050 15.975 3.315 ;
        RECT  11.555 3.085 15.975 3.315 ;
        RECT  15.230 0.970 15.670 1.720 ;
        RECT  15.230 1.380 16.195 1.720 ;
        RECT  13.990 1.540 14.380 1.880 ;
        RECT  14.150 1.540 14.380 2.855 ;
        RECT  15.230 0.970 15.460 2.855 ;
        RECT  14.150 2.570 15.460 2.855 ;
        RECT  14.710 0.410 17.625 0.640 ;
        RECT  12.560 0.970 13.200 1.310 ;
        RECT  14.710 0.410 15.000 1.310 ;
        RECT  12.560 1.080 15.000 1.310 ;
        RECT  17.395 0.410 17.625 1.960 ;
        RECT  17.395 1.620 18.380 1.960 ;
        RECT  12.560 0.970 12.790 2.855 ;
        RECT  12.220 2.515 13.920 2.855 ;
    END
END SDFFSR_X4_18_SVT_WB

MACRO SDFFSR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFSR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.224  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.375 2.270 16.860 3.335 ;
        RECT  16.375 0.870 16.605 3.335 ;
        RECT  16.320 0.870 16.605 1.210 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.960 2.270 18.350 3.280 ;
        RECT  18.025 0.685 18.350 3.280 ;
        RECT  17.960 0.685 18.350 1.440 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.605 1.515 15.100 2.340 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.238  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.010 1.515 13.530 2.155 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 18.480 4.100 ;
        RECT  17.240 2.580 17.580 4.100 ;
        RECT  15.685 3.550 16.025 4.100 ;
        RECT  12.905 3.550 14.455 4.100 ;
        RECT  9.680 3.545 10.020 4.100 ;
        RECT  7.760 3.545 8.100 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 18.480 0.180 ;
        RECT  17.295 -0.180 17.580 1.440 ;
        RECT  14.140 -0.180 14.480 0.825 ;
        RECT  7.940 -0.180 8.280 0.815 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.610 1.100 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  4.430 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.635 1.725 0.870 ;
        RECT  0.470 0.635 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.415 0.930 5.645 3.335 ;
        RECT  2.375 3.105 5.645 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  7.000 2.535 8.680 2.855 ;
        RECT  6.335 0.945 6.685 1.285 ;
        RECT  6.455 1.505 8.900 1.765 ;
        RECT  8.560 1.505 8.900 1.845 ;
        RECT  6.455 0.945 6.685 2.855 ;
        RECT  6.335 2.460 6.685 2.855 ;
        RECT  7.190 1.995 7.530 2.305 ;
        RECT  7.190 2.075 10.185 2.305 ;
        RECT  9.900 0.945 10.185 2.755 ;
        RECT  9.080 2.075 10.185 2.755 ;
        RECT  9.080 2.415 10.725 2.755 ;
        RECT  10.955 1.765 11.345 2.105 ;
        RECT  10.955 1.765 11.185 3.315 ;
        RECT  6.440 3.085 11.185 3.315 ;
        RECT  6.440 3.085 6.780 3.425 ;
        RECT  4.890 0.410 7.255 0.640 ;
        RECT  9.315 0.410 12.320 0.715 ;
        RECT  6.915 0.410 7.255 1.275 ;
        RECT  9.315 0.410 9.655 1.275 ;
        RECT  6.915 1.045 9.655 1.275 ;
        RECT  4.890 0.410 5.120 1.345 ;
        RECT  4.470 1.055 5.120 1.345 ;
        RECT  10.415 0.410 10.665 1.805 ;
        RECT  12.035 0.410 12.320 1.900 ;
        RECT  4.470 1.820 5.040 2.190 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  10.895 0.945 11.180 1.465 ;
        RECT  10.895 1.235 11.805 1.465 ;
        RECT  11.575 1.235 11.805 3.320 ;
        RECT  11.415 2.415 11.805 3.320 ;
        RECT  15.805 2.055 16.145 3.320 ;
        RECT  11.415 3.090 16.145 3.320 ;
        RECT  15.330 0.945 15.670 1.725 ;
        RECT  15.330 1.385 16.145 1.725 ;
        RECT  13.980 1.515 14.375 1.855 ;
        RECT  14.145 1.515 14.375 2.860 ;
        RECT  15.330 0.945 15.560 2.860 ;
        RECT  14.145 2.575 15.560 2.860 ;
        RECT  14.710 0.410 17.065 0.640 ;
        RECT  12.550 0.945 13.290 1.285 ;
        RECT  14.710 0.410 15.050 1.285 ;
        RECT  12.550 1.055 15.050 1.285 ;
        RECT  16.835 0.410 17.065 2.040 ;
        RECT  16.835 1.700 17.795 2.040 ;
        RECT  12.550 0.945 12.780 2.860 ;
        RECT  12.080 2.445 13.900 2.860 ;
    END
END SDFFSR_X2_18_SVT_WB

MACRO SDFFSR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFSR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.224  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.563  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.130 2.790 16.935 3.130 ;
        RECT  16.190 2.290 16.935 3.130 ;
        RECT  16.190 0.980 16.420 3.130 ;
        RECT  16.080 0.980 16.420 1.300 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.400 2.395 17.790 3.365 ;
        RECT  17.510 0.980 17.790 3.365 ;
        RECT  17.400 0.980 17.790 1.320 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.485 1.605 14.980 2.385 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.136  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.238  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.990 1.515 13.510 2.215 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  16.840 3.515 17.170 4.100 ;
        RECT  16.130 3.515 16.425 4.100 ;
        RECT  12.820 3.555 13.730 4.100 ;
        RECT  9.620 3.515 9.960 4.100 ;
        RECT  7.760 3.515 8.100 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  17.110 -0.180 17.450 0.545 ;
        RECT  13.995 -0.180 14.335 0.825 ;
        RECT  8.080 -0.180 8.420 0.815 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.610 1.100 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  4.430 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.635 1.725 0.870 ;
        RECT  0.470 0.635 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.435 0.925 5.665 3.335 ;
        RECT  2.375 3.105 5.665 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  7.000 2.535 8.670 2.825 ;
        RECT  6.335 0.945 6.685 1.285 ;
        RECT  6.455 1.505 8.890 1.735 ;
        RECT  8.550 1.505 8.890 1.835 ;
        RECT  6.455 0.945 6.685 2.825 ;
        RECT  6.335 2.430 6.685 2.825 ;
        RECT  7.190 1.965 7.530 2.305 ;
        RECT  7.190 2.075 10.190 2.305 ;
        RECT  9.890 0.945 10.190 2.750 ;
        RECT  9.085 2.075 10.190 2.750 ;
        RECT  9.085 2.410 10.665 2.750 ;
        RECT  10.895 1.735 11.325 2.075 ;
        RECT  10.895 1.735 11.125 3.285 ;
        RECT  6.440 3.055 11.125 3.285 ;
        RECT  6.440 3.055 6.780 3.385 ;
        RECT  4.890 0.445 7.255 0.675 ;
        RECT  9.320 0.410 12.300 0.715 ;
        RECT  6.915 0.445 7.255 1.275 ;
        RECT  9.320 0.410 9.660 1.275 ;
        RECT  6.915 1.045 9.660 1.275 ;
        RECT  4.890 0.445 5.120 1.375 ;
        RECT  4.470 1.055 5.120 1.375 ;
        RECT  10.420 0.410 10.655 1.805 ;
        RECT  12.015 0.410 12.300 1.855 ;
        RECT  4.470 1.815 5.075 2.195 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  15.210 0.940 15.525 1.910 ;
        RECT  13.845 1.515 14.255 1.840 ;
        RECT  15.210 1.565 15.950 1.910 ;
        RECT  14.025 1.515 14.255 2.865 ;
        RECT  14.025 2.635 15.440 2.865 ;
        RECT  15.210 0.940 15.440 3.045 ;
        RECT  14.700 2.635 15.440 3.045 ;
        RECT  10.885 0.945 11.185 1.455 ;
        RECT  10.885 1.225 11.785 1.455 ;
        RECT  15.670 2.240 15.955 2.580 ;
        RECT  11.555 1.225 11.785 3.325 ;
        RECT  11.355 2.405 11.785 3.325 ;
        RECT  11.355 3.095 14.190 3.325 ;
        RECT  15.670 2.240 15.900 3.505 ;
        RECT  13.955 3.275 15.900 3.505 ;
        RECT  14.640 0.410 16.880 0.710 ;
        RECT  12.530 0.945 13.075 1.285 ;
        RECT  14.640 0.410 14.980 1.285 ;
        RECT  12.530 1.055 14.980 1.285 ;
        RECT  16.650 0.410 16.880 1.935 ;
        RECT  16.650 1.595 17.280 1.935 ;
        RECT  12.530 0.945 12.760 2.785 ;
        RECT  12.020 2.445 13.775 2.785 ;
    END
END SDFFSR_X1_18_SVT_WB

MACRO SDFFSQ_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFSQ_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.505 2.590 16.830 3.405 ;
        RECT  15.035 1.090 16.830 1.360 ;
        RECT  16.505 0.575 16.830 1.360 ;
        RECT  15.035 2.590 16.830 2.925 ;
        RECT  15.705 1.090 16.215 2.925 ;
        RECT  15.035 1.090 16.215 1.365 ;
        RECT  15.035 2.590 15.430 3.410 ;
        RECT  15.035 0.520 15.430 1.365 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.805 1.750 12.195 2.305 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  17.210 3.050 17.550 4.100 ;
        RECT  15.770 3.165 16.110 4.100 ;
        RECT  14.285 3.430 14.635 4.100 ;
        RECT  11.890 3.570 13.170 4.100 ;
        RECT  7.750 3.530 9.030 4.100 ;
        RECT  3.855 3.570 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  17.210 -0.180 17.550 0.815 ;
        RECT  15.770 -0.180 16.110 0.800 ;
        RECT  14.290 -0.180 14.630 0.350 ;
        RECT  12.460 -0.180 12.800 0.350 ;
        RECT  7.600 -0.180 7.940 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.535 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  5.770 0.940 6.120 1.310 ;
        RECT  5.870 0.940 6.120 2.995 ;
        RECT  4.985 2.705 6.120 2.995 ;
        RECT  4.010 1.055 4.240 3.340 ;
        RECT  2.375 3.105 4.240 3.340 ;
        RECT  4.985 2.705 5.215 3.340 ;
        RECT  2.375 3.110 5.215 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.500 1.045 7.080 1.385 ;
        RECT  6.850 2.090 8.460 2.350 ;
        RECT  6.850 1.045 7.080 2.840 ;
        RECT  6.500 2.555 7.080 2.840 ;
        RECT  7.450 1.565 9.075 1.860 ;
        RECT  8.790 1.045 9.075 2.840 ;
        RECT  8.735 1.565 9.075 2.840 ;
        RECT  8.735 2.500 9.910 2.840 ;
        RECT  8.310 2.580 9.910 2.840 ;
        RECT  6.660 3.070 10.080 3.300 ;
        RECT  5.455 3.270 7.100 3.510 ;
        RECT  9.795 3.070 10.080 3.510 ;
        RECT  5.100 0.410 7.100 0.640 ;
        RECT  6.725 0.585 11.110 0.815 ;
        RECT  5.100 0.410 5.330 1.350 ;
        RECT  4.470 1.120 5.330 1.350 ;
        RECT  9.305 0.585 9.535 1.905 ;
        RECT  9.305 1.565 9.620 1.905 ;
        RECT  10.770 0.585 11.110 2.305 ;
        RECT  4.470 2.015 5.525 2.395 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.340 0.865 11.570 2.865 ;
        RECT  11.010 2.580 12.640 2.865 ;
        RECT  9.765 1.045 10.155 1.385 ;
        RECT  10.030 1.180 10.540 1.615 ;
        RECT  13.185 2.005 13.565 2.365 ;
        RECT  10.310 1.180 10.540 3.340 ;
        RECT  10.310 2.530 10.630 3.340 ;
        RECT  13.185 2.005 13.415 3.340 ;
        RECT  10.310 3.105 13.415 3.340 ;
        RECT  12.505 1.045 14.585 1.360 ;
        RECT  12.505 1.045 12.765 1.995 ;
        RECT  14.250 1.640 15.465 1.995 ;
        RECT  14.250 1.045 14.585 2.945 ;
        RECT  13.645 2.595 14.585 2.945 ;
        RECT  13.645 2.595 13.910 3.425 ;
    END
END SDFFSQ_X8_18_SVT_WB

MACRO SDFFSQ_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFSQ_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.035 2.590 16.100 2.925 ;
        RECT  15.780 1.090 16.100 2.925 ;
        RECT  15.035 1.090 16.100 1.365 ;
        RECT  15.035 2.590 15.430 3.410 ;
        RECT  15.035 0.520 15.430 1.365 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.805 1.750 12.195 2.305 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  14.285 3.430 14.635 4.100 ;
        RECT  11.890 3.570 13.170 4.100 ;
        RECT  7.750 3.530 9.030 4.100 ;
        RECT  3.855 3.570 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  14.290 -0.180 14.630 0.350 ;
        RECT  12.460 -0.180 12.800 0.350 ;
        RECT  7.600 -0.180 7.940 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.535 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  5.770 0.940 6.120 1.310 ;
        RECT  5.870 0.940 6.120 2.995 ;
        RECT  4.985 2.705 6.120 2.995 ;
        RECT  4.010 1.055 4.240 3.340 ;
        RECT  2.375 3.105 4.240 3.340 ;
        RECT  4.985 2.705 5.215 3.340 ;
        RECT  2.375 3.110 5.215 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.500 1.045 7.080 1.385 ;
        RECT  6.850 2.090 8.460 2.350 ;
        RECT  6.850 1.045 7.080 2.840 ;
        RECT  6.500 2.555 7.080 2.840 ;
        RECT  7.450 1.565 9.075 1.860 ;
        RECT  8.790 1.045 9.075 2.840 ;
        RECT  8.735 1.565 9.075 2.840 ;
        RECT  8.735 2.500 9.910 2.840 ;
        RECT  8.310 2.580 9.910 2.840 ;
        RECT  6.660 3.070 10.080 3.300 ;
        RECT  5.455 3.270 7.100 3.510 ;
        RECT  9.795 3.070 10.080 3.510 ;
        RECT  5.100 0.410 7.100 0.640 ;
        RECT  6.725 0.585 11.055 0.815 ;
        RECT  5.100 0.410 5.330 1.350 ;
        RECT  4.470 1.120 5.330 1.350 ;
        RECT  9.305 0.585 9.535 1.905 ;
        RECT  9.305 1.565 9.620 1.905 ;
        RECT  10.770 0.585 11.055 2.325 ;
        RECT  4.470 2.015 5.525 2.395 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.305 0.965 11.570 2.875 ;
        RECT  10.990 2.585 12.635 2.875 ;
        RECT  9.765 1.045 10.155 1.385 ;
        RECT  10.030 1.180 10.540 1.615 ;
        RECT  13.185 2.005 13.565 2.365 ;
        RECT  10.310 1.180 10.540 3.340 ;
        RECT  10.310 2.530 10.630 3.340 ;
        RECT  13.185 2.005 13.415 3.340 ;
        RECT  10.310 3.105 13.415 3.340 ;
        RECT  12.505 1.045 14.585 1.360 ;
        RECT  12.505 1.045 12.765 1.995 ;
        RECT  14.250 1.640 15.465 1.995 ;
        RECT  14.250 1.045 14.585 2.945 ;
        RECT  13.645 2.595 14.585 2.945 ;
        RECT  13.645 2.595 13.910 3.425 ;
    END
END SDFFSQ_X4_18_SVT_WB

MACRO SDFFSQ_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFSQ_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.480 2.500 15.545 2.835 ;
        RECT  15.175 1.045 15.545 2.835 ;
        RECT  14.465 1.045 15.545 1.390 ;
        RECT  14.480 2.500 14.865 3.295 ;
        RECT  14.465 0.565 14.785 1.390 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.805 1.750 12.400 2.305 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  12.095 3.570 13.890 4.100 ;
        RECT  7.555 3.530 8.835 4.100 ;
        RECT  3.855 3.570 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  12.665 -0.180 13.975 0.350 ;
        RECT  7.405 -0.180 7.745 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.535 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  5.575 0.940 5.925 1.310 ;
        RECT  5.675 0.940 5.925 2.995 ;
        RECT  4.930 2.705 5.925 2.995 ;
        RECT  4.010 1.055 4.240 3.340 ;
        RECT  2.375 3.105 4.240 3.340 ;
        RECT  4.930 2.705 5.160 3.340 ;
        RECT  2.375 3.110 5.160 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.305 1.045 6.885 1.385 ;
        RECT  6.655 2.090 8.265 2.350 ;
        RECT  6.655 1.045 6.885 2.840 ;
        RECT  6.305 2.555 6.885 2.840 ;
        RECT  7.255 1.565 8.880 1.860 ;
        RECT  8.595 1.045 8.880 2.840 ;
        RECT  8.540 1.565 8.880 2.840 ;
        RECT  8.540 2.500 9.715 2.840 ;
        RECT  8.115 2.580 9.715 2.840 ;
        RECT  6.465 3.070 9.885 3.300 ;
        RECT  5.390 3.270 6.905 3.510 ;
        RECT  9.600 3.070 9.885 3.510 ;
        RECT  5.100 0.410 6.905 0.640 ;
        RECT  6.530 0.585 10.915 0.815 ;
        RECT  5.100 0.410 5.330 1.350 ;
        RECT  4.470 1.055 5.330 1.350 ;
        RECT  9.110 0.585 9.340 1.905 ;
        RECT  9.110 1.565 9.425 1.905 ;
        RECT  4.470 1.055 4.755 2.365 ;
        RECT  10.575 0.585 10.915 2.305 ;
        RECT  4.470 1.985 5.285 2.365 ;
        RECT  4.470 1.055 4.700 2.875 ;
        RECT  11.225 0.910 11.535 2.830 ;
        RECT  10.800 2.575 12.830 2.830 ;
        RECT  9.570 1.045 9.960 1.385 ;
        RECT  9.835 1.180 10.345 1.615 ;
        RECT  13.390 2.005 13.770 2.300 ;
        RECT  10.115 1.180 10.345 3.340 ;
        RECT  10.115 2.530 10.435 3.340 ;
        RECT  13.390 2.005 13.620 3.340 ;
        RECT  10.115 3.105 13.620 3.340 ;
        RECT  12.710 1.045 14.230 1.360 ;
        RECT  12.710 1.045 12.970 1.995 ;
        RECT  14.000 1.645 14.450 1.995 ;
        RECT  14.000 1.045 14.230 2.875 ;
        RECT  13.850 2.530 14.230 2.875 ;
    END
END SDFFSQ_X2_18_SVT_WB

MACRO SDFFSQ_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFSQ_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.480 2.735 15.545 3.070 ;
        RECT  15.175 1.045 15.545 3.070 ;
        RECT  14.465 1.045 15.545 1.390 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.236  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.805 1.750 12.400 2.305 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  15.160 3.515 15.500 4.100 ;
        RECT  12.095 3.570 13.375 4.100 ;
        RECT  7.555 3.530 8.835 4.100 ;
        RECT  3.855 3.570 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  15.160 -0.180 15.500 0.405 ;
        RECT  12.665 -0.180 13.005 0.350 ;
        RECT  7.405 -0.180 7.745 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.535 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.185 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.185 0.580 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  5.575 0.940 5.925 1.310 ;
        RECT  5.675 0.940 5.925 2.995 ;
        RECT  4.930 2.705 5.925 2.995 ;
        RECT  4.010 1.055 4.240 3.340 ;
        RECT  2.375 3.105 4.240 3.340 ;
        RECT  4.930 2.705 5.160 3.340 ;
        RECT  2.375 3.110 5.160 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.305 1.045 6.885 1.385 ;
        RECT  6.655 2.090 8.265 2.350 ;
        RECT  6.655 1.045 6.885 2.840 ;
        RECT  6.305 2.555 6.885 2.840 ;
        RECT  7.255 1.565 8.880 1.860 ;
        RECT  8.595 1.045 8.880 2.840 ;
        RECT  8.540 1.565 8.880 2.840 ;
        RECT  8.540 2.500 9.715 2.840 ;
        RECT  8.115 2.580 9.715 2.840 ;
        RECT  6.465 3.070 9.885 3.300 ;
        RECT  5.390 3.270 6.905 3.510 ;
        RECT  9.600 3.070 9.885 3.510 ;
        RECT  5.100 0.410 6.905 0.640 ;
        RECT  6.530 0.585 10.915 0.815 ;
        RECT  5.100 0.410 5.330 1.350 ;
        RECT  4.470 1.055 5.330 1.350 ;
        RECT  9.110 0.585 9.340 1.905 ;
        RECT  9.110 1.565 9.425 1.905 ;
        RECT  4.470 1.055 4.755 2.365 ;
        RECT  10.575 0.585 10.915 2.305 ;
        RECT  4.470 1.985 5.285 2.365 ;
        RECT  4.470 1.055 4.700 2.875 ;
        RECT  11.185 0.970 11.505 2.845 ;
        RECT  10.795 2.570 12.825 2.845 ;
        RECT  9.570 1.045 9.960 1.385 ;
        RECT  9.835 1.180 10.345 1.615 ;
        RECT  13.390 2.005 13.770 2.300 ;
        RECT  10.115 1.180 10.345 3.340 ;
        RECT  10.115 2.530 10.435 3.340 ;
        RECT  13.390 2.005 13.620 3.340 ;
        RECT  10.115 3.105 13.620 3.340 ;
        RECT  12.710 1.100 14.230 1.360 ;
        RECT  12.710 1.100 12.970 1.995 ;
        RECT  14.000 1.645 14.450 1.995 ;
        RECT  14.000 1.100 14.230 2.875 ;
        RECT  13.850 2.530 14.230 2.875 ;
    END
END SDFFSQ_X1_18_SVT_WB

MACRO SDFFR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.135 1.100 14.460 3.310 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.605 0.540 16.170 3.385 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.275  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.920 3.250 12.365 3.510 ;
        RECT  8.920 1.920 9.150 3.510 ;
        RECT  6.860 1.920 9.150 2.170 ;
        RECT  6.860 1.770 7.285 2.170 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.800 4.100 ;
        RECT  14.845 3.045 15.185 4.100 ;
        RECT  12.825 3.515 13.655 4.100 ;
        RECT  8.405 3.050 8.690 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.800 0.180 ;
        RECT  14.845 -0.180 15.185 0.405 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.560 1.040 1.915 1.335 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  5.350 0.875 5.645 1.225 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.195 2.435 5.580 3.340 ;
        RECT  2.375 3.105 4.705 3.335 ;
        RECT  5.350 0.875 5.580 3.340 ;
        RECT  4.540 3.110 5.580 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.800 2.400 8.405 2.740 ;
        RECT  6.025 0.875 7.735 1.215 ;
        RECT  7.505 0.875 7.735 1.690 ;
        RECT  7.505 1.445 9.145 1.690 ;
        RECT  6.340 0.875 6.570 2.770 ;
        RECT  5.935 2.430 6.570 2.770 ;
        RECT  7.965 0.875 9.610 1.215 ;
        RECT  9.380 0.875 9.610 3.020 ;
        RECT  4.890 0.410 10.530 0.645 ;
        RECT  4.890 0.410 5.120 1.340 ;
        RECT  4.470 1.055 5.120 1.340 ;
        RECT  10.300 0.410 10.530 2.500 ;
        RECT  4.470 1.815 5.065 2.190 ;
        RECT  10.300 2.160 10.550 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.755 1.465 12.845 1.805 ;
        RECT  9.840 0.875 10.070 3.020 ;
        RECT  11.755 1.465 12.035 3.020 ;
        RECT  9.840 2.730 12.035 3.020 ;
        RECT  11.240 0.875 13.305 1.215 ;
        RECT  13.075 0.875 13.305 3.015 ;
        RECT  11.240 0.875 11.525 1.860 ;
        RECT  13.075 1.860 13.460 3.015 ;
        RECT  12.265 2.675 13.460 3.015 ;
        RECT  10.760 0.415 14.455 0.645 ;
        RECT  13.885 0.635 15.375 0.870 ;
        RECT  10.760 0.415 11.010 1.215 ;
        RECT  15.035 0.635 15.375 1.960 ;
        RECT  10.780 0.415 11.010 2.500 ;
        RECT  10.780 2.160 11.175 2.500 ;
    END
END SDFFR_X4_18_SVT_WB

MACRO SDFFR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.885 1.100 14.300 2.765 ;
        RECT  13.575 2.375 13.910 3.310 ;
        RECT  13.575 1.100 14.300 1.455 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.100 0.540 15.540 3.385 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.275  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.920 3.250 12.365 3.510 ;
        RECT  8.920 1.920 9.150 3.510 ;
        RECT  6.860 1.920 9.150 2.170 ;
        RECT  6.860 1.770 7.285 2.170 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  14.285 3.045 14.625 4.100 ;
        RECT  12.825 3.515 13.180 4.100 ;
        RECT  8.405 3.050 8.690 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  14.285 -0.180 14.625 0.405 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.560 1.040 1.915 1.335 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  5.350 0.875 5.645 1.225 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.195 2.435 5.580 3.340 ;
        RECT  2.375 3.105 4.705 3.335 ;
        RECT  5.350 0.875 5.580 3.340 ;
        RECT  4.540 3.110 5.580 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.800 2.400 8.405 2.740 ;
        RECT  6.025 0.875 7.735 1.215 ;
        RECT  7.505 0.875 7.735 1.690 ;
        RECT  7.505 1.445 9.145 1.690 ;
        RECT  6.340 0.875 6.570 2.770 ;
        RECT  5.935 2.430 6.570 2.770 ;
        RECT  7.965 0.875 9.610 1.215 ;
        RECT  9.380 0.875 9.610 3.020 ;
        RECT  4.890 0.410 10.530 0.645 ;
        RECT  4.890 0.410 5.120 1.340 ;
        RECT  4.470 1.055 5.120 1.340 ;
        RECT  10.300 0.410 10.530 2.500 ;
        RECT  4.470 1.815 5.065 2.190 ;
        RECT  10.300 2.160 10.550 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.755 1.465 12.845 1.805 ;
        RECT  9.840 0.875 10.070 3.020 ;
        RECT  11.755 1.465 12.035 3.020 ;
        RECT  9.840 2.730 12.035 3.020 ;
        RECT  11.240 0.875 13.305 1.215 ;
        RECT  11.240 0.875 11.525 1.860 ;
        RECT  13.075 1.910 13.545 2.145 ;
        RECT  13.075 0.875 13.305 3.015 ;
        RECT  12.265 2.675 13.305 3.015 ;
        RECT  10.760 0.415 13.895 0.645 ;
        RECT  13.595 0.635 14.815 0.870 ;
        RECT  10.760 0.415 11.010 1.215 ;
        RECT  14.530 0.635 14.815 1.975 ;
        RECT  10.780 0.415 11.010 2.500 ;
        RECT  10.780 2.160 11.175 2.500 ;
    END
END SDFFR_X2_18_SVT_WB

MACRO SDFFR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.885 1.100 14.300 2.765 ;
        RECT  13.575 2.375 13.910 3.405 ;
        RECT  13.575 1.100 14.300 1.455 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.100 1.075 15.540 3.385 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.275  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.920 3.250 12.365 3.510 ;
        RECT  8.920 1.920 9.150 3.510 ;
        RECT  6.860 1.920 9.150 2.170 ;
        RECT  6.860 1.770 7.285 2.170 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  14.285 3.045 14.625 4.100 ;
        RECT  12.825 3.515 13.180 4.100 ;
        RECT  8.405 3.050 8.690 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  14.285 -0.180 14.625 0.405 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.560 1.040 1.915 1.335 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  5.350 0.875 5.645 1.225 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.195 2.435 5.580 3.340 ;
        RECT  2.375 3.105 4.705 3.335 ;
        RECT  5.350 0.875 5.580 3.340 ;
        RECT  4.540 3.110 5.580 3.340 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.800 2.400 8.405 2.740 ;
        RECT  6.025 0.875 7.735 1.215 ;
        RECT  7.505 0.875 7.735 1.690 ;
        RECT  7.505 1.445 9.145 1.690 ;
        RECT  6.340 0.875 6.570 2.770 ;
        RECT  5.935 2.430 6.570 2.770 ;
        RECT  7.965 0.875 9.610 1.215 ;
        RECT  9.380 0.875 9.610 3.020 ;
        RECT  4.890 0.410 10.530 0.645 ;
        RECT  4.890 0.410 5.120 1.340 ;
        RECT  4.470 1.055 5.120 1.340 ;
        RECT  10.300 0.410 10.530 2.500 ;
        RECT  4.470 1.815 5.065 2.190 ;
        RECT  10.300 2.160 10.550 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.755 1.465 12.845 1.805 ;
        RECT  9.840 0.875 10.070 3.020 ;
        RECT  11.755 1.465 12.035 3.020 ;
        RECT  9.840 2.730 12.035 3.020 ;
        RECT  11.240 0.875 13.305 1.215 ;
        RECT  11.240 0.875 11.525 1.860 ;
        RECT  13.075 1.910 13.545 2.145 ;
        RECT  13.075 0.875 13.305 3.015 ;
        RECT  12.265 2.675 13.305 3.015 ;
        RECT  10.760 0.415 13.895 0.645 ;
        RECT  13.595 0.635 14.815 0.870 ;
        RECT  10.760 0.415 11.010 1.215 ;
        RECT  14.530 0.635 14.815 1.975 ;
        RECT  10.780 0.415 11.010 2.500 ;
        RECT  10.780 2.160 11.175 2.500 ;
    END
END SDFFR_X1_18_SVT_WB

MACRO SDFFRQ_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFRQ_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.300  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.785 0.535 15.125 3.450 ;
        RECT  13.465 1.620 15.125 1.955 ;
        RECT  13.465 0.540 13.885 3.450 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.030 3.250 12.080 3.510 ;
        RECT  9.030 1.920 9.260 3.510 ;
        RECT  6.860 1.920 9.260 2.150 ;
        RECT  6.860 1.770 7.370 2.150 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  15.505 2.625 15.845 4.100 ;
        RECT  12.745 3.165 13.085 4.100 ;
        RECT  8.515 3.050 8.800 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  15.505 -0.180 15.845 1.440 ;
        RECT  12.705 -0.180 13.045 0.405 ;
        RECT  11.000 -0.180 11.340 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.545 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.465 0.410 4.700 0.825 ;
        RECT  3.245 0.595 4.700 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.415 0.875 5.645 3.335 ;
        RECT  2.375 3.105 5.645 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.855 2.380 8.500 2.720 ;
        RECT  6.855 2.380 7.140 3.000 ;
        RECT  6.080 0.875 7.870 1.215 ;
        RECT  7.590 0.875 7.870 1.690 ;
        RECT  7.590 1.445 9.245 1.690 ;
        RECT  6.395 0.875 6.625 2.720 ;
        RECT  6.080 2.380 6.625 2.720 ;
        RECT  8.100 0.875 9.725 1.215 ;
        RECT  9.490 0.875 9.725 3.020 ;
        RECT  4.955 0.410 10.645 0.645 ;
        RECT  4.955 0.410 5.185 1.345 ;
        RECT  4.470 1.055 5.185 1.345 ;
        RECT  10.415 0.410 10.645 2.500 ;
        RECT  4.470 1.790 5.140 2.220 ;
        RECT  10.415 2.160 10.785 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.410 1.860 12.540 2.200 ;
        RECT  9.955 0.875 10.185 3.020 ;
        RECT  11.410 1.860 11.750 3.020 ;
        RECT  9.955 2.730 11.750 3.020 ;
        RECT  12.205 0.875 12.545 1.630 ;
        RECT  10.875 1.395 13.230 1.630 ;
        RECT  10.875 1.395 11.205 1.735 ;
        RECT  12.890 1.395 13.230 2.935 ;
        RECT  11.980 2.625 13.230 2.935 ;
    END
END SDFFRQ_X8_18_SVT_WB

MACRO SDFFRQ_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFRQ_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.465 0.540 13.885 3.450 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.030 3.250 12.080 3.510 ;
        RECT  9.030 1.920 9.260 3.510 ;
        RECT  6.860 1.920 9.260 2.150 ;
        RECT  6.860 1.770 7.370 2.150 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.560 4.100 ;
        RECT  12.745 3.165 13.085 4.100 ;
        RECT  8.515 3.050 8.800 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.560 0.180 ;
        RECT  12.705 -0.180 13.045 0.405 ;
        RECT  11.000 -0.180 11.340 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.545 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.465 0.410 4.700 0.825 ;
        RECT  3.245 0.595 4.700 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.415 0.875 5.645 3.335 ;
        RECT  2.375 3.105 5.645 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.855 2.380 8.500 2.720 ;
        RECT  6.855 2.380 7.140 3.000 ;
        RECT  6.080 0.875 7.870 1.215 ;
        RECT  7.590 0.875 7.870 1.690 ;
        RECT  7.590 1.445 9.245 1.690 ;
        RECT  6.395 0.875 6.625 2.720 ;
        RECT  6.080 2.380 6.625 2.720 ;
        RECT  8.100 0.875 9.725 1.215 ;
        RECT  9.490 0.875 9.725 3.020 ;
        RECT  4.955 0.410 10.645 0.645 ;
        RECT  4.955 0.410 5.185 1.345 ;
        RECT  4.470 1.055 5.185 1.345 ;
        RECT  10.415 0.410 10.645 2.500 ;
        RECT  4.470 1.790 5.140 2.220 ;
        RECT  10.415 2.160 10.785 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.410 1.860 12.540 2.200 ;
        RECT  9.955 0.875 10.185 3.020 ;
        RECT  11.410 1.860 11.750 3.020 ;
        RECT  9.955 2.730 11.750 3.020 ;
        RECT  12.205 0.875 12.545 1.630 ;
        RECT  10.875 1.395 13.230 1.630 ;
        RECT  10.875 1.395 11.205 1.735 ;
        RECT  12.890 1.395 13.230 2.935 ;
        RECT  11.980 2.625 13.230 2.935 ;
    END
END SDFFRQ_X4_18_SVT_WB

MACRO SDFFRQ_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFRQ_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.465 0.540 13.860 3.450 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.030 3.250 12.080 3.510 ;
        RECT  9.030 1.920 9.260 3.510 ;
        RECT  6.860 1.920 9.260 2.150 ;
        RECT  6.860 1.770 7.370 2.150 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.000 4.100 ;
        RECT  12.745 3.165 13.085 4.100 ;
        RECT  8.515 3.050 8.800 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.000 0.180 ;
        RECT  12.705 -0.180 13.045 0.405 ;
        RECT  11.000 -0.180 11.340 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.545 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.465 0.410 4.700 0.825 ;
        RECT  3.245 0.595 4.700 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.415 0.875 5.645 3.335 ;
        RECT  2.375 3.105 5.645 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.855 2.380 8.500 2.720 ;
        RECT  6.855 2.380 7.140 3.000 ;
        RECT  6.080 0.875 7.870 1.215 ;
        RECT  7.590 0.875 7.870 1.690 ;
        RECT  7.590 1.445 9.245 1.690 ;
        RECT  6.395 0.875 6.625 2.720 ;
        RECT  6.080 2.380 6.625 2.720 ;
        RECT  8.100 0.875 9.725 1.215 ;
        RECT  9.490 0.875 9.725 3.020 ;
        RECT  4.955 0.410 10.645 0.645 ;
        RECT  4.955 0.410 5.185 1.345 ;
        RECT  4.470 1.055 5.185 1.345 ;
        RECT  10.415 0.410 10.645 2.500 ;
        RECT  4.470 1.790 5.140 2.220 ;
        RECT  10.415 2.160 10.785 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.410 1.860 12.540 2.200 ;
        RECT  9.955 0.875 10.185 3.020 ;
        RECT  11.410 1.860 11.750 3.020 ;
        RECT  9.955 2.730 11.750 3.020 ;
        RECT  12.205 0.875 12.545 1.630 ;
        RECT  10.875 1.395 13.230 1.630 ;
        RECT  10.875 1.395 11.205 1.735 ;
        RECT  12.890 1.395 13.230 2.935 ;
        RECT  11.980 2.625 13.230 2.935 ;
    END
END SDFFRQ_X2_18_SVT_WB

MACRO SDFFRQ_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFRQ_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.465 0.540 13.860 3.450 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.191  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.030 3.250 12.080 3.510 ;
        RECT  9.030 1.920 9.260 3.510 ;
        RECT  6.860 1.920 9.260 2.150 ;
        RECT  6.860 1.770 7.370 2.150 ;
        END
    END RN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.000 4.100 ;
        RECT  12.745 3.165 13.085 4.100 ;
        RECT  8.515 3.050 8.800 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.000 0.180 ;
        RECT  12.705 -0.180 13.045 0.405 ;
        RECT  11.000 -0.180 11.340 0.355 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.545 1.040 1.915 1.325 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.465 0.410 4.700 0.825 ;
        RECT  3.245 0.595 4.700 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.415 0.875 5.645 3.335 ;
        RECT  2.375 3.105 5.645 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.855 2.380 8.500 2.720 ;
        RECT  6.855 2.380 7.140 3.000 ;
        RECT  6.080 0.875 7.870 1.215 ;
        RECT  7.590 0.875 7.870 1.690 ;
        RECT  7.590 1.445 9.245 1.690 ;
        RECT  6.395 0.875 6.625 2.720 ;
        RECT  6.080 2.380 6.625 2.720 ;
        RECT  8.100 0.875 9.725 1.215 ;
        RECT  9.490 0.875 9.725 3.020 ;
        RECT  4.955 0.410 10.645 0.645 ;
        RECT  4.955 0.410 5.185 1.345 ;
        RECT  4.470 1.055 5.185 1.345 ;
        RECT  10.415 0.410 10.645 2.500 ;
        RECT  4.470 1.790 5.140 2.220 ;
        RECT  10.415 2.160 10.785 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  11.410 1.860 12.540 2.200 ;
        RECT  9.955 0.875 10.185 3.020 ;
        RECT  11.410 1.860 11.750 3.020 ;
        RECT  9.955 2.730 11.750 3.020 ;
        RECT  12.205 0.875 12.545 1.630 ;
        RECT  10.875 1.395 13.230 1.630 ;
        RECT  10.875 1.395 11.205 1.735 ;
        RECT  12.890 1.395 13.230 2.935 ;
        RECT  11.980 2.625 13.230 2.935 ;
    END
END SDFFRQ_X1_18_SVT_WB

MACRO SDFFQ_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFQ_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.300  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.120 0.540 13.460 3.330 ;
        RECT  11.800 1.615 13.460 1.950 ;
        RECT  11.800 0.535 12.190 3.325 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.560 4.100 ;
        RECT  13.840 2.385 14.190 4.100 ;
        RECT  9.975 3.515 11.385 4.100 ;
        RECT  7.265 2.705 7.605 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.560 0.180 ;
        RECT  13.840 -0.180 14.180 1.395 ;
        RECT  11.040 -0.180 11.380 0.405 ;
        RECT  9.780 -0.180 10.120 0.410 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.540 1.040 1.915 1.330 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.350 0.880 5.580 3.335 ;
        RECT  2.375 3.105 5.580 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.575 1.220 ;
        RECT  7.345 0.880 7.575 1.740 ;
        RECT  7.345 1.400 7.775 1.740 ;
        RECT  6.290 0.880 6.520 2.995 ;
        RECT  6.015 2.655 6.520 2.995 ;
        RECT  7.805 0.880 8.325 1.170 ;
        RECT  6.750 1.990 7.025 2.475 ;
        RECT  6.750 2.135 8.325 2.475 ;
        RECT  8.005 0.880 8.325 3.020 ;
        RECT  7.985 2.135 8.325 3.020 ;
        RECT  4.890 0.410 9.370 0.650 ;
        RECT  4.890 0.410 5.120 1.340 ;
        RECT  4.470 1.055 5.120 1.340 ;
        RECT  4.470 1.820 5.025 2.240 ;
        RECT  9.070 0.410 9.370 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.650 2.085 10.660 2.425 ;
        RECT  8.555 0.880 8.840 3.020 ;
        RECT  9.650 2.085 9.990 3.020 ;
        RECT  8.555 2.730 9.990 3.020 ;
        RECT  10.540 0.880 10.880 1.830 ;
        RECT  9.600 1.490 10.880 1.830 ;
        RECT  9.600 1.600 11.350 1.830 ;
        RECT  11.010 1.600 11.350 3.015 ;
        RECT  10.540 2.675 11.350 3.015 ;
    END
END SDFFQ_X8_18_SVT_WB

MACRO SDFFQ_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFQ_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.800 0.535 12.190 3.325 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  9.975 3.515 11.385 4.100 ;
        RECT  7.265 2.705 7.605 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  11.040 -0.180 11.380 0.405 ;
        RECT  9.780 -0.180 10.120 0.410 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.540 1.040 1.915 1.330 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.350 0.880 5.580 3.335 ;
        RECT  2.375 3.105 5.580 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.575 1.220 ;
        RECT  7.345 0.880 7.575 1.740 ;
        RECT  7.345 1.400 7.775 1.740 ;
        RECT  6.290 0.880 6.520 2.995 ;
        RECT  6.015 2.655 6.520 2.995 ;
        RECT  7.805 0.880 8.325 1.170 ;
        RECT  6.750 1.990 7.025 2.475 ;
        RECT  6.750 2.135 8.325 2.475 ;
        RECT  8.005 0.880 8.325 3.020 ;
        RECT  7.985 2.135 8.325 3.020 ;
        RECT  4.890 0.410 9.370 0.650 ;
        RECT  4.890 0.410 5.120 1.340 ;
        RECT  4.470 1.055 5.120 1.340 ;
        RECT  4.470 1.820 5.025 2.240 ;
        RECT  9.070 0.410 9.370 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.650 2.085 10.660 2.425 ;
        RECT  8.555 0.880 8.840 3.020 ;
        RECT  9.650 2.085 9.990 3.020 ;
        RECT  8.555 2.730 9.990 3.020 ;
        RECT  10.540 0.880 10.880 1.830 ;
        RECT  9.600 1.490 10.880 1.830 ;
        RECT  9.600 1.600 11.350 1.830 ;
        RECT  11.010 1.600 11.350 3.015 ;
        RECT  10.540 2.675 11.350 3.015 ;
    END
END SDFFQ_X4_18_SVT_WB

MACRO SDFFQ_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFQ_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.800 0.535 12.180 3.325 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  9.975 3.515 11.385 4.100 ;
        RECT  7.265 2.705 7.605 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.040 -0.180 11.380 0.405 ;
        RECT  9.780 -0.180 10.120 0.410 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.540 1.040 1.915 1.330 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.350 0.880 5.580 3.335 ;
        RECT  2.375 3.105 5.580 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.575 1.220 ;
        RECT  7.345 0.880 7.575 1.740 ;
        RECT  7.345 1.400 7.775 1.740 ;
        RECT  6.290 0.880 6.520 2.995 ;
        RECT  6.015 2.655 6.520 2.995 ;
        RECT  7.805 0.880 8.325 1.170 ;
        RECT  6.750 1.990 7.025 2.475 ;
        RECT  6.750 2.135 8.325 2.475 ;
        RECT  8.005 0.880 8.325 3.020 ;
        RECT  7.985 2.135 8.325 3.020 ;
        RECT  4.890 0.410 9.370 0.650 ;
        RECT  4.890 0.410 5.120 1.340 ;
        RECT  4.470 1.055 5.120 1.340 ;
        RECT  4.470 1.820 5.025 2.240 ;
        RECT  9.070 0.410 9.370 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.650 2.085 10.660 2.425 ;
        RECT  8.555 0.880 8.840 3.020 ;
        RECT  9.650 2.085 9.990 3.020 ;
        RECT  8.555 2.730 9.990 3.020 ;
        RECT  10.540 0.880 10.880 1.830 ;
        RECT  9.600 1.490 10.880 1.830 ;
        RECT  9.600 1.600 11.350 1.830 ;
        RECT  11.010 1.600 11.350 3.015 ;
        RECT  10.540 2.675 11.350 3.015 ;
    END
END SDFFQ_X2_18_SVT_WB

MACRO SDFFQ_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFQ_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.800 0.535 12.180 3.325 ;
        END
    END Q
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  9.975 3.515 11.385 4.100 ;
        RECT  7.265 2.705 7.605 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.040 -0.180 11.380 0.405 ;
        RECT  9.780 -0.180 10.120 0.410 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.540 1.040 1.915 1.330 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.350 0.880 5.580 3.335 ;
        RECT  2.375 3.105 5.580 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.575 1.220 ;
        RECT  7.345 0.880 7.575 1.740 ;
        RECT  7.345 1.400 7.775 1.740 ;
        RECT  6.290 0.880 6.520 2.995 ;
        RECT  6.015 2.655 6.520 2.995 ;
        RECT  7.805 0.880 8.325 1.170 ;
        RECT  6.750 1.990 7.025 2.475 ;
        RECT  6.750 2.135 8.325 2.475 ;
        RECT  8.005 0.880 8.325 3.020 ;
        RECT  7.985 2.135 8.325 3.020 ;
        RECT  4.890 0.410 9.370 0.650 ;
        RECT  4.890 0.410 5.120 1.340 ;
        RECT  4.470 1.055 5.120 1.340 ;
        RECT  4.470 1.820 5.025 2.240 ;
        RECT  9.070 0.410 9.370 2.500 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.650 2.085 10.660 2.425 ;
        RECT  8.555 0.880 8.840 3.020 ;
        RECT  9.650 2.085 9.990 3.020 ;
        RECT  8.555 2.730 9.990 3.020 ;
        RECT  10.540 0.880 10.880 1.830 ;
        RECT  9.600 1.490 10.880 1.830 ;
        RECT  9.600 1.600 11.350 1.830 ;
        RECT  11.010 1.600 11.350 3.015 ;
        RECT  10.540 2.675 11.350 3.015 ;
    END
END SDFFQ_X1_18_SVT_WB

MACRO SDFFQN_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFQN_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.800 0.590 12.215 3.450 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  9.950 3.455 11.350 4.100 ;
        RECT  7.280 2.650 7.620 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  11.040 -0.180 11.380 0.460 ;
        RECT  9.780 -0.180 10.120 0.445 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.560 1.040 1.915 1.330 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.350 0.880 5.580 3.335 ;
        RECT  2.375 3.105 5.580 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.580 1.220 ;
        RECT  7.350 0.880 7.580 1.740 ;
        RECT  7.350 1.400 7.805 1.740 ;
        RECT  6.335 0.880 6.565 2.985 ;
        RECT  6.020 2.645 6.565 2.985 ;
        RECT  7.810 0.880 8.285 1.170 ;
        RECT  6.795 1.955 7.025 2.420 ;
        RECT  6.795 2.080 8.285 2.420 ;
        RECT  8.035 0.880 8.285 2.985 ;
        RECT  8.000 2.080 8.285 2.985 ;
        RECT  4.890 0.410 9.330 0.650 ;
        RECT  4.890 0.410 5.120 1.350 ;
        RECT  4.470 1.055 5.120 1.350 ;
        RECT  4.470 1.835 5.115 2.180 ;
        RECT  9.045 0.410 9.330 2.465 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.845 1.915 10.640 2.145 ;
        RECT  8.530 0.880 8.815 2.985 ;
        RECT  9.845 1.915 10.075 2.985 ;
        RECT  8.530 2.695 10.075 2.985 ;
        RECT  10.540 0.880 10.880 1.685 ;
        RECT  9.560 1.400 11.100 1.685 ;
        RECT  10.870 1.400 11.100 2.980 ;
        RECT  10.540 2.640 11.100 2.980 ;
    END
END SDFFQN_X4_18_SVT_WB

MACRO SDFFQN_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFQN_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.800 0.590 12.180 3.450 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  9.950 3.455 11.350 4.100 ;
        RECT  7.280 2.650 7.620 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.040 -0.180 11.380 0.460 ;
        RECT  9.780 -0.180 10.120 0.445 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.560 1.040 1.915 1.330 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.350 0.880 5.580 3.335 ;
        RECT  2.375 3.105 5.580 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.580 1.220 ;
        RECT  7.350 0.880 7.580 1.740 ;
        RECT  7.350 1.400 7.805 1.740 ;
        RECT  6.335 0.880 6.565 2.985 ;
        RECT  6.020 2.645 6.565 2.985 ;
        RECT  7.810 0.880 8.285 1.170 ;
        RECT  6.795 1.955 7.025 2.420 ;
        RECT  6.795 2.080 8.285 2.420 ;
        RECT  8.035 0.880 8.285 2.985 ;
        RECT  8.000 2.080 8.285 2.985 ;
        RECT  4.890 0.410 9.330 0.650 ;
        RECT  4.890 0.410 5.120 1.350 ;
        RECT  4.470 1.055 5.120 1.350 ;
        RECT  4.470 1.835 5.115 2.180 ;
        RECT  9.045 0.410 9.330 2.465 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.845 1.915 10.640 2.145 ;
        RECT  8.530 0.880 8.815 2.985 ;
        RECT  9.845 1.915 10.075 2.985 ;
        RECT  8.530 2.695 10.075 2.985 ;
        RECT  10.540 0.880 10.880 1.685 ;
        RECT  9.560 1.400 11.100 1.685 ;
        RECT  10.870 1.400 11.100 2.980 ;
        RECT  10.540 2.640 11.100 2.980 ;
    END
END SDFFQN_X2_18_SVT_WB

MACRO SDFFQN_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN SDFFQN_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.102  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.245 3.085 0.980 3.315 ;
        RECT  0.700 2.855 0.980 3.315 ;
        RECT  0.245 3.085 0.585 3.510 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.245  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.770 3.780 2.150 ;
        RECT  2.890 1.515 3.400 1.800 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.800 0.590 12.180 3.450 ;
        END
    END QN
    PIN SE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.620 1.380 1.960 ;
        RECT  0.700 1.620 1.040 2.190 ;
        END
    END SE
    PIN SI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.115  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 2.130 2.940 2.415 ;
        RECT  2.145 1.770 2.660 2.415 ;
        RECT  2.145 0.990 2.485 2.415 ;
        END
    END SI
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  9.950 3.455 11.350 4.100 ;
        RECT  7.280 2.650 7.620 4.100 ;
        RECT  3.855 3.565 4.195 4.100 ;
        RECT  0.815 3.545 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.040 -0.180 11.380 0.460 ;
        RECT  9.780 -0.180 10.120 0.445 ;
        RECT  3.855 -0.180 4.195 0.365 ;
        RECT  0.815 -0.180 1.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.560 1.040 1.915 1.330 ;
        RECT  1.610 1.040 1.915 2.875 ;
        RECT  3.335 2.535 3.675 2.875 ;
        RECT  1.610 2.645 3.675 2.875 ;
        RECT  1.385 0.410 3.585 0.660 ;
        RECT  0.470 0.580 1.725 0.810 ;
        RECT  4.425 0.410 4.660 0.825 ;
        RECT  3.245 0.595 4.660 0.825 ;
        RECT  0.470 0.580 0.810 1.160 ;
        RECT  0.185 0.930 0.470 2.855 ;
        RECT  2.715 0.890 3.005 1.285 ;
        RECT  2.715 1.055 4.240 1.285 ;
        RECT  4.010 1.055 4.240 3.335 ;
        RECT  5.350 0.880 5.580 3.335 ;
        RECT  2.375 3.105 5.580 3.335 ;
        RECT  2.375 3.105 2.715 3.420 ;
        RECT  6.015 0.880 7.580 1.220 ;
        RECT  7.350 0.880 7.580 1.740 ;
        RECT  7.350 1.400 7.805 1.740 ;
        RECT  6.335 0.880 6.565 2.985 ;
        RECT  6.020 2.645 6.565 2.985 ;
        RECT  7.810 0.880 8.285 1.170 ;
        RECT  6.795 1.955 7.025 2.420 ;
        RECT  6.795 2.080 8.285 2.420 ;
        RECT  8.035 0.880 8.285 2.985 ;
        RECT  8.000 2.080 8.285 2.985 ;
        RECT  4.890 0.410 9.330 0.650 ;
        RECT  4.890 0.410 5.120 1.350 ;
        RECT  4.470 1.055 5.120 1.350 ;
        RECT  4.470 1.835 5.115 2.180 ;
        RECT  9.045 0.410 9.330 2.465 ;
        RECT  4.470 1.055 4.755 2.875 ;
        RECT  9.845 1.915 10.640 2.145 ;
        RECT  8.530 0.880 8.815 2.985 ;
        RECT  9.845 1.915 10.075 2.985 ;
        RECT  8.530 2.695 10.075 2.985 ;
        RECT  10.540 0.880 10.880 1.685 ;
        RECT  9.560 1.400 11.100 1.685 ;
        RECT  10.870 1.400 11.100 2.980 ;
        RECT  10.540 2.640 11.100 2.980 ;
    END
END SDFFQN_X1_18_SVT_WB

MACRO OR4_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR4_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 2.240 3.630 2.470 ;
        RECT  2.820 1.915 3.630 2.470 ;
        RECT  1.810 2.240 2.150 2.715 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.000 1.455 4.340 2.150 ;
        RECT  2.120 1.455 4.340 1.685 ;
        RECT  2.120 1.455 2.460 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.620 0.995 5.045 1.920 ;
        RECT  1.470 0.995 5.045 1.225 ;
        RECT  1.470 0.995 1.770 1.960 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.670 2.150 5.775 2.380 ;
        RECT  5.435 1.900 5.775 2.380 ;
        RECT  2.380 2.700 4.990 2.930 ;
        RECT  4.670 2.150 4.990 2.930 ;
        RECT  0.735 2.945 2.720 3.285 ;
        RECT  2.380 2.700 2.720 3.285 ;
        RECT  0.735 1.840 1.020 3.285 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.456  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.115 0.685 8.455 1.440 ;
        RECT  7.980 2.640 8.390 3.270 ;
        RECT  8.025 1.440 8.390 3.270 ;
        RECT  6.670 1.440 8.390 1.670 ;
        RECT  6.490 2.640 8.390 2.870 ;
        RECT  6.670 0.685 7.010 1.670 ;
        RECT  6.490 2.640 6.830 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  8.835 2.545 9.175 4.100 ;
        RECT  7.290 3.100 7.630 4.100 ;
        RECT  5.730 3.070 6.070 4.100 ;
        RECT  0.180 2.615 0.505 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  8.835 -0.180 9.175 1.375 ;
        RECT  7.395 -0.180 7.735 1.210 ;
        RECT  5.950 -0.180 6.290 1.210 ;
        RECT  0.180 -0.180 0.520 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.470 5.560 0.765 ;
        RECT  0.900 0.470 1.240 1.225 ;
        RECT  5.275 0.470 5.560 1.670 ;
        RECT  5.275 1.440 6.260 1.670 ;
        RECT  6.030 1.900 7.410 2.200 ;
        RECT  6.030 1.440 6.260 2.840 ;
        RECT  5.220 2.610 6.260 2.840 ;
        RECT  5.220 2.610 5.500 3.450 ;
        RECT  3.060 3.160 5.500 3.450 ;
    END
END OR4_X8_18_SVT_WB

MACRO OR4_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR4_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.640 0.670 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.380 1.490 2.720 ;
        RECT  1.150 1.860 1.490 2.720 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 2.390 2.380 2.730 ;
        RECT  1.810 1.860 2.150 2.730 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.670 2.905 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.080 1.850 5.420 3.385 ;
        RECT  3.675 1.060 5.420 1.400 ;
        RECT  5.080 0.590 5.420 1.400 ;
        RECT  3.675 1.850 5.420 2.190 ;
        RECT  4.560 1.060 4.900 2.190 ;
        RECT  3.675 1.850 3.980 3.385 ;
        RECT  3.675 0.535 3.980 1.400 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.360 2.575 4.700 4.100 ;
        RECT  2.880 3.515 3.220 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.360 -0.180 4.700 0.810 ;
        RECT  2.880 -0.180 3.220 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.800 0.630 1.140 1.440 ;
        RECT  2.120 0.535 2.460 1.440 ;
        RECT  0.800 1.100 2.460 1.440 ;
        RECT  0.800 1.105 3.445 1.440 ;
        RECT  3.160 1.105 3.445 3.285 ;
        RECT  0.240 3.055 3.445 3.285 ;
        RECT  0.240 3.055 0.580 3.450 ;
    END
END OR4_X6_18_SVT_WB

MACRO OR4_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR4_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.595 1.760 1.090 2.175 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.440 1.260 1.780 1.960 ;
        RECT  1.210 1.260 1.780 1.550 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.110 1.260 2.845 1.600 ;
        RECT  2.110 1.260 2.450 1.960 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.790 1.910 3.220 2.710 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.257  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.000 0.535 4.340 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.720 2.580 5.060 4.100 ;
        RECT  3.180 3.515 3.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.720 -0.180 5.060 1.345 ;
        RECT  3.240 -0.180 3.580 0.405 ;
        RECT  1.720 -0.180 2.060 0.405 ;
        RECT  0.240 -0.180 0.580 1.390 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.480 0.535 2.820 0.920 ;
        RECT  0.960 0.635 3.770 0.920 ;
        RECT  0.530 2.405 0.870 3.280 ;
        RECT  3.460 0.635 3.770 3.280 ;
        RECT  0.530 2.940 3.770 3.280 ;
    END
END OR4_X4_18_SVT_WB

MACRO OR4_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR4_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.440 0.940 2.770 ;
        RECT  0.140 2.320 0.445 2.770 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.580 1.540 2.180 ;
        RECT  0.960 1.580 1.540 1.985 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.630 2.310 2.105 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.125 2.335 2.725 2.780 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.415 2.590 3.780 3.270 ;
        RECT  3.500 0.535 3.780 3.270 ;
        RECT  3.415 0.535 3.780 1.445 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  2.640 3.515 2.980 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.925 -0.180 2.960 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.040 3.185 1.280 ;
        RECT  2.955 1.850 3.270 2.200 ;
        RECT  2.955 1.040 3.185 3.240 ;
        RECT  0.330 3.010 3.185 3.240 ;
    END
END OR4_X2_18_SVT_WB

MACRO OR4_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR4_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.755 0.795 2.150 ;
        RECT  0.450 1.615 0.795 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.435 1.585 1.785 ;
        RECT  1.260 1.080 1.585 1.785 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.580 2.035 2.100 2.370 ;
        RECT  1.815 1.595 2.100 2.370 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.162  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.480 2.660 2.290 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 2.260 3.780 2.990 ;
        RECT  3.550 0.670 3.780 2.990 ;
        RECT  3.420 0.670 3.780 1.015 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  2.625 3.515 2.965 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.185 -0.180 0.490 0.480 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.745 0.475 2.405 0.705 ;
        RECT  2.055 0.475 2.405 1.060 ;
        RECT  2.055 0.830 3.190 1.060 ;
        RECT  0.745 0.475 1.030 1.205 ;
        RECT  2.905 1.315 3.320 1.620 ;
        RECT  2.905 0.830 3.190 2.925 ;
        RECT  0.245 2.635 3.190 2.925 ;
    END
END OR4_X1_18_SVT_WB

MACRO OR4_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR4_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 2.140 3.550 2.370 ;
        RECT  2.740 1.915 3.550 2.370 ;
        RECT  1.820 2.140 2.160 2.710 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.455 4.340 2.150 ;
        RECT  2.040 1.455 4.340 1.685 ;
        RECT  2.040 1.455 2.380 1.910 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.610 0.995 4.950 1.980 ;
        RECT  1.405 0.995 4.950 1.225 ;
        RECT  1.405 0.995 1.670 1.960 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.390 2.600 5.630 2.830 ;
        RECT  5.320 1.860 5.630 2.830 ;
        RECT  0.945 2.940 2.730 3.280 ;
        RECT  2.390 2.600 2.730 3.280 ;
        RECT  0.945 1.760 1.175 3.280 ;
        RECT  0.460 1.760 1.175 2.180 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.360 0.590 9.700 3.330 ;
        RECT  8.080 1.520 9.700 1.860 ;
        RECT  7.840 2.380 8.310 3.330 ;
        RECT  8.080 1.520 8.310 3.330 ;
        RECT  6.400 1.440 8.260 1.670 ;
        RECT  7.840 0.590 8.260 1.670 ;
        RECT  6.320 2.380 8.310 2.720 ;
        RECT  6.400 0.590 6.740 1.670 ;
        RECT  6.320 2.380 6.660 3.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  10.080 2.630 10.480 4.100 ;
        RECT  8.600 2.630 8.940 4.100 ;
        RECT  7.040 3.100 7.435 4.100 ;
        RECT  5.560 3.520 5.900 4.100 ;
        RECT  0.180 2.470 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  10.080 -0.180 10.475 1.290 ;
        RECT  8.600 -0.180 8.940 1.290 ;
        RECT  7.120 -0.180 7.460 1.210 ;
        RECT  0.180 -0.180 0.520 1.375 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.470 6.090 0.755 ;
        RECT  5.860 1.900 7.850 2.150 ;
        RECT  5.860 0.470 6.090 3.290 ;
        RECT  2.980 3.060 6.090 3.290 ;
        RECT  2.980 3.060 3.320 3.400 ;
    END
END OR4_X12_18_SVT_WB

MACRO OR3_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR3_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.040 1.820 2.710 2.180 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.130 1.620 3.640 1.960 ;
        RECT  3.130 1.260 3.360 1.960 ;
        RECT  1.220 1.260 3.360 1.590 ;
        RECT  1.220 1.260 1.560 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.580 2.410 4.390 2.660 ;
        RECT  4.010 1.840 4.390 2.660 ;
        RECT  0.580 1.860 0.890 2.660 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.660 0.525 7.000 3.395 ;
        RECT  5.220 2.250 7.000 2.480 ;
        RECT  6.250 1.040 7.000 2.480 ;
        RECT  5.220 1.040 7.000 1.280 ;
        RECT  5.220 2.250 5.560 3.190 ;
        RECT  5.220 0.525 5.560 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.940 2.710 6.280 4.100 ;
        RECT  4.460 3.515 4.800 4.100 ;
        RECT  0.310 3.045 0.650 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.940 -0.180 6.280 0.810 ;
        RECT  4.500 -0.180 4.840 0.740 ;
        RECT  3.020 -0.180 3.360 0.350 ;
        RECT  1.500 -0.180 1.840 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.580 4.120 0.875 ;
        RECT  3.780 0.580 4.120 1.200 ;
        RECT  3.780 0.970 4.990 1.200 ;
        RECT  4.760 1.620 5.735 1.960 ;
        RECT  4.760 0.970 4.990 3.285 ;
        RECT  2.260 2.945 4.990 3.285 ;
    END
END OR3_X8_18_SVT_WB

MACRO OR3_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR3_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.940 1.210 2.320 1.695 ;
        RECT  1.635 1.210 2.320 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.925 3.645 2.165 ;
        RECT  2.860 1.755 3.645 2.165 ;
        RECT  1.240 1.825 1.560 2.165 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.780 2.395 4.340 2.625 ;
        RECT  4.000 1.445 4.340 2.625 ;
        RECT  0.780 1.820 1.010 2.625 ;
        RECT  0.465 1.820 1.010 2.160 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.660 2.495 7.000 3.385 ;
        RECT  5.220 0.990 7.000 1.255 ;
        RECT  6.660 0.470 7.000 1.255 ;
        RECT  5.220 2.495 7.000 2.830 ;
        RECT  5.730 0.990 6.130 2.830 ;
        RECT  5.220 2.495 5.560 3.385 ;
        RECT  5.220 0.470 5.560 1.255 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.940 3.100 6.280 4.100 ;
        RECT  4.460 3.515 4.800 4.100 ;
        RECT  0.310 2.825 0.650 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  5.940 -0.180 6.280 0.760 ;
        RECT  4.500 -0.180 4.840 0.755 ;
        RECT  3.020 -0.180 3.360 0.405 ;
        RECT  1.500 -0.180 1.840 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.635 4.120 0.975 ;
        RECT  3.780 0.635 4.120 1.215 ;
        RECT  3.780 0.985 4.990 1.215 ;
        RECT  4.705 1.745 5.390 2.040 ;
        RECT  4.705 0.985 4.990 3.160 ;
        RECT  2.260 2.855 4.990 3.160 ;
    END
END OR3_X6_18_SVT_WB

MACRO OR3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.820 1.175 2.180 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.405 1.260 1.745 1.960 ;
        RECT  1.175 1.260 1.745 1.590 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.360 2.415 2.700 ;
        RECT  2.075 1.840 2.415 2.700 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.205  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.260 1.770 3.830 2.135 ;
        RECT  3.260 0.980 3.560 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.940 2.580 4.280 4.100 ;
        RECT  2.445 3.515 2.785 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.940 -0.180 4.280 1.280 ;
        RECT  2.460 -0.180 2.800 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 0.635 3.030 0.975 ;
        RECT  0.170 0.635 0.520 1.455 ;
        RECT  0.495 2.410 0.835 3.270 ;
        RECT  2.745 0.635 3.030 3.270 ;
        RECT  0.495 2.930 3.030 3.270 ;
    END
END OR3_X4_18_SVT_WB

MACRO OR3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.330 1.000 2.775 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.730 1.470 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.625 2.140 2.160 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 2.380 3.220 3.385 ;
        RECT  2.990 0.580 3.220 3.385 ;
        RECT  2.840 0.580 3.220 1.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.080 3.515 2.420 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.035 -0.180 2.390 0.410 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.055 2.610 1.395 ;
        RECT  2.380 1.620 2.760 1.960 ;
        RECT  1.615 2.875 2.610 3.215 ;
        RECT  2.380 1.055 2.610 3.215 ;
        RECT  0.460 3.075 1.800 3.415 ;
    END
END OR3_X2_18_SVT_WB

MACRO OR3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 2.155 1.080 2.480 ;
        RECT  0.115 1.770 0.420 2.480 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.485 1.540 1.825 ;
        RECT  0.650 1.260 1.030 1.825 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.485 2.185 2.100 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.875 0.860 3.220 3.075 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.080 3.515 2.420 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.040 -0.180 2.385 0.405 ;
        RECT  0.940 -0.180 1.280 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.550 0.520 1.030 ;
        RECT  0.180 0.800 2.645 1.030 ;
        RECT  1.500 0.800 2.645 1.255 ;
        RECT  2.415 0.800 2.645 2.940 ;
        RECT  0.540 2.710 2.645 2.940 ;
        RECT  0.540 2.710 0.880 3.050 ;
    END
END OR3_X1_18_SVT_WB

MACRO OR3_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR3_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.660 1.090 2.180 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.980 1.455 5.320 1.905 ;
        RECT  3.600 1.455 5.320 1.685 ;
        RECT  2.840 1.760 3.870 2.100 ;
        RECT  3.600 1.455 3.870 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.100 2.135 6.630 2.365 ;
        RECT  6.180 1.820 6.630 2.365 ;
        RECT  4.100 1.915 4.440 2.365 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.020 2.570 10.360 3.390 ;
        RECT  7.380 0.950 10.360 1.280 ;
        RECT  10.020 0.470 10.360 1.280 ;
        RECT  7.380 2.570 10.360 2.900 ;
        RECT  8.700 2.570 9.040 3.390 ;
        RECT  8.700 0.470 9.040 1.280 ;
        RECT  8.495 0.950 8.885 2.900 ;
        RECT  7.380 2.570 7.720 3.390 ;
        RECT  7.380 0.470 7.720 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  6.660 3.110 7.000 4.100 ;
        RECT  3.820 3.525 4.160 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  6.660 -0.180 7.000 0.810 ;
        RECT  5.220 -0.180 5.560 0.755 ;
        RECT  3.780 -0.180 4.120 0.755 ;
        RECT  2.340 -0.180 2.680 0.755 ;
        RECT  0.900 -0.180 1.240 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 3.065 5.560 3.295 ;
        RECT  5.220 3.065 5.560 3.450 ;
        RECT  0.180 0.670 0.520 1.225 ;
        RECT  0.180 0.985 6.280 1.225 ;
        RECT  5.940 1.040 7.150 1.325 ;
        RECT  6.865 1.690 8.035 1.980 ;
        RECT  6.865 1.040 7.150 2.825 ;
        RECT  0.180 2.595 7.150 2.825 ;
        RECT  0.180 2.595 0.520 3.405 ;
    END
END OR3_X12_18_SVT_WB

MACRO OR2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.710 1.620 2.280 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.500 2.330 2.840 2.660 ;
        RECT  2.510 1.840 2.840 2.660 ;
        RECT  0.500 1.620 0.840 2.660 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.020 2.485 5.360 3.385 ;
        RECT  3.580 1.040 5.360 1.370 ;
        RECT  5.020 0.470 5.360 1.370 ;
        RECT  3.580 2.485 5.360 2.800 ;
        RECT  4.535 1.040 4.925 2.800 ;
        RECT  3.580 2.485 3.920 3.385 ;
        RECT  3.580 0.535 3.920 1.370 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.300 3.095 4.640 4.100 ;
        RECT  0.310 3.110 0.650 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.300 -0.180 4.640 0.810 ;
        RECT  1.500 -0.180 1.840 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.535 1.080 1.345 ;
        RECT  2.260 0.535 2.600 1.345 ;
        RECT  0.740 1.105 3.350 1.345 ;
        RECT  3.120 1.630 3.760 1.965 ;
        RECT  3.120 1.105 3.350 3.220 ;
        RECT  1.540 2.890 3.350 3.220 ;
    END
END OR2_X8_18_SVT_WB

MACRO OR2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.245 1.195 1.850 1.720 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.950 2.750 2.180 ;
        RECT  2.410 1.840 2.750 2.180 ;
        RECT  0.140 1.770 0.790 2.180 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.050 2.510 5.390 3.385 ;
        RECT  3.610 0.990 5.390 1.290 ;
        RECT  5.050 0.470 5.390 1.290 ;
        RECT  3.610 2.510 5.390 2.795 ;
        RECT  4.600 0.990 4.950 2.795 ;
        RECT  3.610 2.510 3.950 3.385 ;
        RECT  3.610 0.470 3.950 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.330 3.095 4.670 4.100 ;
        RECT  2.850 3.515 3.190 4.100 ;
        RECT  0.300 2.820 0.640 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.330 -0.180 4.670 0.760 ;
        RECT  2.890 -0.180 3.230 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.725 0.690 2.510 0.965 ;
        RECT  2.170 0.690 2.510 1.215 ;
        RECT  0.725 0.690 1.070 1.030 ;
        RECT  2.170 0.985 3.380 1.215 ;
        RECT  3.095 1.630 3.805 1.970 ;
        RECT  3.095 0.985 3.380 2.750 ;
        RECT  1.450 2.410 3.380 2.750 ;
    END
END OR2_X6_18_SVT_WB

MACRO OR2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.580 0.665 1.960 ;
        RECT  0.140 1.160 0.470 1.960 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.615 2.340 1.375 2.710 ;
        RECT  1.090 1.840 1.375 2.710 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.075 2.575 3.220 2.915 ;
        RECT  2.905 1.055 3.220 2.915 ;
        RECT  2.075 1.055 3.220 1.355 ;
        RECT  2.075 2.575 2.455 3.385 ;
        RECT  2.075 0.535 2.455 1.355 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.790 3.165 3.130 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.780 -0.180 3.120 0.805 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.755 0.690 1.835 1.030 ;
        RECT  1.605 1.650 2.235 1.920 ;
        RECT  1.605 0.690 1.835 3.280 ;
        RECT  0.180 2.940 1.835 3.280 ;
    END
END OR2_X4_18_SVT_WB

MACRO OR2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.105 0.760 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.820 1.405 2.175 ;
        RECT  1.020 1.575 1.405 2.175 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.095 2.580 2.660 3.390 ;
        RECT  2.340 0.470 2.660 3.390 ;
        RECT  2.245 0.470 2.660 1.325 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  1.330 3.105 1.670 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.180 -0.180 0.520 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.470 1.925 0.810 ;
        RECT  1.635 0.470 1.925 2.135 ;
        RECT  1.635 1.765 2.110 2.135 ;
        RECT  1.635 0.470 1.865 2.875 ;
        RECT  0.180 2.645 1.865 2.875 ;
        RECT  0.180 2.645 0.520 3.295 ;
    END
END OR2_X2_18_SVT_WB

MACRO OR2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.205 0.980 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.205 1.590 1.835 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.540 2.660 3.380 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  1.520 3.100 1.860 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.220 -0.180 0.480 0.985 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.645 2.050 0.975 ;
        RECT  1.820 0.645 2.050 2.870 ;
        RECT  0.330 2.640 2.050 2.870 ;
        RECT  0.330 2.640 0.670 3.225 ;
    END
END OR2_X1_18_SVT_WB

MACRO OR2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN OR2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.540 1.455 2.880 1.905 ;
        RECT  0.915 1.455 2.880 1.685 ;
        RECT  0.395 1.805 1.255 2.200 ;
        RECT  0.915 1.455 1.255 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.485 2.135 4.080 2.365 ;
        RECT  3.445 1.750 4.080 2.365 ;
        RECT  1.485 1.915 1.845 2.365 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.820 2.495 8.160 3.390 ;
        RECT  4.940 0.990 8.160 1.275 ;
        RECT  7.820 0.470 8.160 1.275 ;
        RECT  4.940 2.495 8.160 2.800 ;
        RECT  6.380 0.985 8.160 1.275 ;
        RECT  6.380 2.495 6.720 3.390 ;
        RECT  6.380 0.470 6.720 1.275 ;
        RECT  6.290 0.990 6.630 2.800 ;
        RECT  4.940 2.495 5.280 3.390 ;
        RECT  4.940 0.470 5.280 1.275 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  7.100 3.150 7.440 4.100 ;
        RECT  5.660 3.150 6.000 4.100 ;
        RECT  4.220 3.110 4.560 4.100 ;
        RECT  1.340 3.110 1.680 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  7.100 -0.180 7.440 0.755 ;
        RECT  5.660 -0.180 6.000 0.760 ;
        RECT  4.220 -0.180 4.560 0.765 ;
        RECT  2.780 -0.180 3.120 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.520 1.080 1.225 ;
        RECT  2.050 0.485 2.410 1.225 ;
        RECT  3.490 0.455 3.835 1.225 ;
        RECT  0.740 0.995 4.710 1.225 ;
        RECT  4.425 1.650 6.015 2.005 ;
        RECT  4.425 0.995 4.710 2.880 ;
        RECT  0.180 2.595 4.710 2.880 ;
        RECT  0.180 2.595 0.520 3.405 ;
        RECT  2.780 2.595 3.120 3.405 ;
    END
END OR2_X12_18_SVT_WB

MACRO OAI33_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI33_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.770 1.760 3.220 2.215 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.485 1.620 3.830 2.210 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.620 4.535 2.205 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.760 2.405 3.220 ;
        RECT  2.100 1.620 2.405 3.220 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.230 1.620 1.740 2.150 ;
        RECT  1.230 1.620 1.460 2.475 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.535 1.745 1.000 2.180 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.655 0.470 7.140 2.885 ;
        RECT  6.655 0.470 6.980 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.920 2.695 6.260 4.100 ;
        RECT  4.490 3.045 4.830 4.100 ;
        RECT  0.430 2.460 0.770 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.920 -0.180 6.260 0.810 ;
        RECT  1.620 -0.180 1.960 0.905 ;
        RECT  0.180 -0.180 0.520 1.320 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.340 0.565 4.120 0.860 ;
        RECT  0.900 1.035 1.240 1.375 ;
        RECT  2.340 0.565 2.680 1.375 ;
        RECT  0.900 1.135 2.680 1.375 ;
        RECT  4.500 0.620 4.840 1.375 ;
        RECT  3.060 1.090 4.995 1.375 ;
        RECT  4.765 1.775 5.780 2.005 ;
        RECT  4.765 1.010 4.995 2.785 ;
        RECT  2.635 2.445 4.995 2.785 ;
        RECT  2.635 2.445 2.920 3.255 ;
        RECT  5.225 0.565 5.540 1.545 ;
        RECT  5.225 1.315 6.425 1.545 ;
        RECT  6.165 1.315 6.425 2.465 ;
        RECT  5.225 2.235 6.425 2.465 ;
        RECT  5.225 2.235 5.540 3.215 ;
    END
END OAI33_X4_18_SVT_WB

MACRO OAI33_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI33_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.760 1.760 3.220 2.205 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.620 3.800 2.320 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.620 4.395 2.320 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.660 2.440 1.960 ;
        RECT  1.770 2.380 2.300 2.765 ;
        RECT  2.070 1.660 2.300 2.765 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.660 1.720 2.100 ;
        RECT  1.210 1.660 1.440 2.330 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.515 1.745 0.980 2.180 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.910  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.530 2.550 4.910 2.785 ;
        RECT  4.625 0.650 4.910 2.785 ;
        RECT  3.060 1.155 4.910 1.390 ;
        RECT  4.500 0.650 4.910 1.390 ;
        RECT  2.530 2.445 2.870 3.255 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.390 3.015 4.730 4.100 ;
        RECT  0.430 2.460 0.770 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.620 -0.180 1.960 0.970 ;
        RECT  0.180 -0.180 0.520 1.385 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.340 0.630 4.120 0.925 ;
        RECT  0.900 1.100 1.240 1.430 ;
        RECT  2.340 0.630 2.680 1.430 ;
        RECT  0.900 1.200 2.680 1.430 ;
    END
END OAI33_X2_18_SVT_WB

MACRO OAI33_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI33_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.375 2.330 2.875 2.830 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.640 3.500 2.100 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 2.330 4.155 2.830 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.580 2.180 2.145 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.375 1.660 3.035 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.785 1.030 2.230 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.846  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 3.060 4.900 3.305 ;
        RECT  4.620 1.045 4.900 3.305 ;
        RECT  2.890 1.045 4.900 1.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.380 3.535 4.720 4.100 ;
        RECT  0.310 2.990 0.650 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.500 -0.180 1.840 1.340 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
END OAI33_X1_18_SVT_WB

MACRO OAI33_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI33_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.565 1.260 2.905 2.000 ;
        RECT  2.330 1.260 2.905 1.540 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.305 2.305 3.780 2.710 ;
        RECT  3.305 1.950 3.645 2.710 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.055 1.620 4.340 2.430 ;
        RECT  3.875 1.620 4.340 2.075 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.815 1.740 2.215 2.245 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.250 2.465 1.740 3.270 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.950 1.020 2.760 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 2.940 4.860 3.230 ;
        RECT  4.570 0.560 4.860 3.230 ;
        RECT  3.135 1.030 4.860 1.370 ;
        RECT  4.520 0.560 4.860 1.370 ;
        RECT  3.135 1.030 3.420 1.540 ;
        RECT  2.330 2.940 2.700 3.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.270 3.460 4.610 4.100 ;
        RECT  0.445 2.995 0.830 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.640 -0.180 1.980 1.440 ;
        RECT  0.180 -0.180 0.520 0.875 ;
        END
    END VSS
END OAI33_X0_18_SVT_WB

MACRO OAI32_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI32_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.985 1.645 2.710 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.330 3.550 2.690 ;
        RECT  3.170 1.820 3.550 2.690 ;
        RECT  1.260 1.860 1.600 2.690 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.990 1.095 4.330 2.060 ;
        RECT  0.520 1.095 4.330 1.415 ;
        RECT  0.130 1.640 0.860 2.200 ;
        RECT  0.520 1.095 0.860 2.200 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.595 2.240 6.245 2.745 ;
        RECT  5.865 1.915 6.245 2.745 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.745 1.455 7.215 2.130 ;
        RECT  5.020 1.455 7.215 1.685 ;
        RECT  5.020 1.455 5.305 2.060 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.560 0.995 6.935 1.225 ;
        RECT  5.875 3.055 6.215 3.450 ;
        RECT  2.220 3.055 6.215 3.285 ;
        RECT  2.220 2.940 4.790 3.285 ;
        RECT  4.560 0.995 4.790 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  7.025 2.640 7.365 4.100 ;
        RECT  4.325 3.515 4.665 4.100 ;
        RECT  0.180 2.640 0.480 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  2.255 -0.180 2.605 0.370 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.980 0.495 7.655 0.765 ;
        RECT  0.180 0.600 4.250 0.865 ;
        RECT  7.315 0.495 7.655 1.230 ;
    END
END OAI32_X4_18_SVT_WB

MACRO OAI32_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI32_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.210 2.190 1.960 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.630 1.585 2.185 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.770 0.980 2.190 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.655 3.270 2.355 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.770 4.070 2.175 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.464  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.105 3.520 1.425 ;
        RECT  2.380 2.890 2.800 3.340 ;
        RECT  2.430 2.585 2.800 3.340 ;
        RECT  2.430 1.105 2.660 3.340 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.900 2.445 4.240 4.100 ;
        RECT  0.220 2.460 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  1.700 -0.180 2.040 0.405 ;
        RECT  0.220 -0.180 0.560 1.385 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.460 0.535 2.800 0.875 ;
        RECT  0.940 0.635 4.240 0.875 ;
        RECT  0.940 0.635 1.280 1.360 ;
        RECT  3.900 0.635 4.240 1.385 ;
    END
END OAI32_X2_18_SVT_WB

MACRO OAI32_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI32_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.615 2.170 2.100 ;
        RECT  1.720 1.615 2.050 2.250 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 2.925 1.610 3.220 ;
        RECT  1.270 2.915 1.610 3.220 ;
        RECT  1.270 2.410 1.505 3.220 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.335 2.335 1.040 2.695 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 2.330 2.770 2.850 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.460 2.390 3.780 3.270 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.000 0.965 3.290 1.570 ;
        RECT  2.115 3.080 3.230 3.335 ;
        RECT  3.000 0.965 3.230 3.335 ;
        RECT  2.810 0.965 3.290 1.565 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.395 3.565 3.740 4.100 ;
        RECT  0.180 3.045 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.500 -0.180 1.840 1.375 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
END OAI32_X1_18_SVT_WB

MACRO OAI32_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI32_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.600 1.635 2.115 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.030 2.880 1.600 3.220 ;
        RECT  1.260 2.525 1.600 3.220 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.220 0.710 2.815 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.770 2.700 2.445 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.390 2.250 3.780 2.865 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.200 2.875 3.160 3.105 ;
        RECT  2.930 1.065 3.160 3.105 ;
        RECT  2.840 1.065 3.160 1.405 ;
        RECT  2.200 2.875 2.660 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.390 3.095 3.730 4.100 ;
        RECT  0.180 3.045 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.500 -0.180 1.840 1.405 ;
        RECT  0.180 -0.180 0.520 0.865 ;
        END
    END VSS
END OAI32_X0_18_SVT_WB

MACRO OAI31_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI31_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.770 2.950 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.180 1.150 3.520 2.060 ;
        RECT  1.810 1.150 3.520 1.540 ;
        RECT  1.190 1.740 2.040 2.080 ;
        RECT  1.810 1.150 2.040 2.080 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.731  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.795 1.765 4.135 2.060 ;
        RECT  0.300 2.380 4.055 2.660 ;
        RECT  3.795 1.765 4.055 2.660 ;
        RECT  0.300 1.860 0.640 2.660 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.535 2.140 5.125 2.710 ;
        RECT  4.535 1.860 4.825 2.710 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.814  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.085 2.940 5.775 3.280 ;
        RECT  5.495 1.090 5.775 3.280 ;
        RECT  4.835 1.090 5.775 1.405 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.490 3.560 5.835 4.100 ;
        RECT  0.180 3.110 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  0.720 -0.180 1.085 0.415 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.350 0.580 5.925 0.845 ;
        RECT  4.140 0.580 4.480 1.295 ;
        RECT  1.350 0.580 1.580 1.305 ;
        RECT  0.180 1.060 1.580 1.305 ;
    END
END OAI31_X4_18_SVT_WB

MACRO OAI31_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI31_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.610 2.495 2.370 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.340 1.590 2.660 ;
        RECT  1.290 1.625 1.590 2.660 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.655 1.035 2.185 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.770 1.510 3.220 2.330 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.167  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.635 2.560 3.780 2.815 ;
        RECT  3.450 0.630 3.780 2.815 ;
        RECT  2.635 2.560 2.975 3.370 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.395 3.045 3.735 4.100 ;
        RECT  0.395 2.435 0.735 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.875 -0.180 2.215 0.820 ;
        RECT  0.395 -0.180 0.735 1.385 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.635 0.470 2.975 1.280 ;
        RECT  1.115 1.050 2.975 1.280 ;
        RECT  1.115 0.620 1.455 1.395 ;
    END
END OAI31_X2_18_SVT_WB

MACRO OAI31_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI31_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.890 2.045 3.230 ;
        RECT  1.760 2.040 2.045 3.230 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.320 1.430 2.660 ;
        RECT  1.090 2.040 1.430 2.660 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.210 0.800 1.590 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.770 2.780 2.340 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.325 2.575 3.240 2.925 ;
        RECT  3.010 0.625 3.240 2.925 ;
        RECT  2.840 0.625 3.240 1.030 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.220 3.460 2.975 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.520 -0.180 1.860 1.350 ;
        RECT  0.180 -0.180 0.520 0.965 ;
        END
    END VSS
END OAI31_X1_18_SVT_WB

MACRO OAI31_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI31_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.580 2.150 2.105 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.330 1.600 2.940 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 2.245 1.020 2.865 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.305 2.780 2.680 ;
        RECT  2.440 2.145 2.780 2.680 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 3.045 3.240 3.385 ;
        RECT  3.010 1.065 3.240 3.385 ;
        RECT  2.840 1.065 3.240 1.590 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.275 3.100 0.690 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.500 -0.180 1.840 1.350 ;
        RECT  0.180 -0.180 0.520 0.865 ;
        END
    END VSS
END OAI31_X0_18_SVT_WB

MACRO OAI22_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI22_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.250 2.880 2.765 3.220 ;
        RECT  2.250 1.640 2.535 3.220 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.745 3.270 2.280 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.260 1.515 1.960 ;
        RECT  0.650 1.260 1.515 1.600 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.140 0.890 2.370 ;
        RECT  0.550 1.860 0.890 2.370 ;
        RECT  0.140 2.140 0.540 2.710 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.160 0.525 7.500 3.395 ;
        RECT  5.720 2.640 7.500 2.980 ;
        RECT  7.125 0.940 7.500 2.980 ;
        RECT  5.720 0.940 7.500 1.280 ;
        RECT  5.720 2.640 6.060 3.395 ;
        RECT  5.720 0.525 6.060 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.880 2.420 8.220 4.100 ;
        RECT  4.960 3.515 5.300 4.100 ;
        RECT  3.180 2.740 3.520 4.100 ;
        RECT  0.270 2.990 0.610 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.880 -0.180 8.220 1.280 ;
        RECT  4.960 -0.180 5.300 0.405 ;
        RECT  0.940 -0.180 1.280 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.580 3.480 0.875 ;
        RECT  1.745 1.105 4.220 1.410 ;
        RECT  3.990 1.105 4.220 2.010 ;
        RECT  3.990 1.670 4.915 2.010 ;
        RECT  1.745 1.105 2.020 3.190 ;
        RECT  4.450 1.100 5.375 1.440 ;
        RECT  5.145 1.620 6.705 1.960 ;
        RECT  5.145 1.100 5.375 2.720 ;
        RECT  4.400 2.380 5.375 2.720 ;
    END
END OAI22_X8_18_SVT_WB

MACRO OAI22_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI22_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.530 1.915 5.340 2.660 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.630 1.760 6.070 2.100 ;
        RECT  5.630 1.455 5.970 2.100 ;
        RECT  4.060 1.455 5.970 1.685 ;
        RECT  3.820 1.685 4.300 1.980 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.560 1.770 2.370 2.265 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.260 3.130 1.960 ;
        RECT  0.870 1.260 3.130 1.540 ;
        RECT  0.870 1.260 1.175 2.200 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.600 0.995 5.820 1.225 ;
        RECT  1.800 2.945 5.100 3.285 ;
        RECT  3.360 1.225 3.830 1.455 ;
        RECT  1.800 2.940 3.590 3.285 ;
        RECT  3.360 1.225 3.590 3.285 ;
        RECT  1.800 2.495 2.140 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  5.920 2.435 6.260 4.100 ;
        RECT  3.280 3.515 3.620 4.100 ;
        RECT  0.180 2.490 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  2.560 -0.180 2.900 0.405 ;
        RECT  0.980 -0.180 1.320 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.170 0.470 6.540 0.765 ;
        RECT  0.220 0.635 3.370 0.975 ;
        RECT  6.200 0.470 6.540 1.225 ;
        RECT  0.220 0.470 0.560 1.280 ;
    END
END OAI22_X4_18_SVT_WB

MACRO OAI22_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI22_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.640 2.670 2.975 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.690 3.440 2.310 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.300 1.260 1.590 1.960 ;
        RECT  1.115 1.260 1.590 1.540 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.165 1.735 0.980 2.315 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.130 2.845 1.410 ;
        RECT  1.820 1.130 2.100 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.225 2.615 3.565 4.100 ;
        RECT  0.395 2.615 0.735 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.975 -0.180 1.315 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.215 0.635 3.565 0.900 ;
        RECT  3.225 0.635 3.565 1.360 ;
        RECT  0.215 0.635 0.555 1.400 ;
    END
END OAI22_X2_18_SVT_WB

MACRO OAI22_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI22_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.400 2.365 2.160 2.785 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 2.375 3.220 3.270 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.115 1.510 1.620 2.115 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.435 2.345 1.030 2.770 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.390 0.925 2.735 1.630 ;
        RECT  1.685 3.100 2.620 3.330 ;
        RECT  2.390 0.925 2.620 3.330 ;
        RECT  2.270 0.925 2.735 1.625 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.350 3.045 0.695 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.790 -0.180 1.140 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.235 1.030 1.895 1.260 ;
    END
END OAI22_X1_18_SVT_WB

MACRO OAI22_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI22_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.660 2.365 2.150 2.785 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 2.000 3.220 2.810 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.555 1.430 2.260 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.490 0.725 2.815 ;
        RECT  0.130 1.920 0.470 2.815 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.575 3.015 2.660 3.330 ;
        RECT  2.380 0.985 2.660 3.330 ;
        RECT  2.245 0.985 2.660 1.325 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.425 3.045 0.765 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.295 -0.180 1.105 0.585 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.985 1.865 1.325 ;
    END
END OAI22_X0_18_SVT_WB

MACRO OAI222_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI222_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.950 1.620 9.315 1.960 ;
        RECT  7.180 1.455 9.290 1.685 ;
        RECT  6.860 1.620 7.410 1.960 ;
        RECT  6.860 1.620 7.175 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.890 1.915 8.700 2.660 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 1.455 6.540 1.960 ;
        RECT  3.570 1.455 6.540 1.685 ;
        RECT  3.570 1.455 4.390 2.100 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.000 1.915 5.810 2.660 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.455 3.220 2.180 ;
        RECT  0.750 1.455 3.220 1.685 ;
        RECT  0.750 1.455 1.060 1.960 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.430 1.915 2.240 2.660 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.296  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.545 0.995 9.775 2.940 ;
        RECT  0.500 2.940 9.610 3.285 ;
        RECT  9.270 2.585 9.775 2.940 ;
        RECT  7.400 0.995 9.775 1.225 ;
        RECT  6.680 2.515 7.020 3.285 ;
        RECT  0.500 2.505 0.840 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  8.080 3.515 8.420 4.100 ;
        RECT  5.200 3.515 5.540 4.100 ;
        RECT  1.700 3.515 2.040 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  3.100 -0.180 3.440 0.765 ;
        RECT  1.660 -0.180 2.000 0.765 ;
        RECT  0.180 -0.180 0.520 0.995 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.525 1.280 1.225 ;
        RECT  2.380 0.525 2.720 1.225 ;
        RECT  0.940 0.995 6.300 1.225 ;
        RECT  3.800 0.470 9.900 0.765 ;
        RECT  6.680 0.470 7.020 1.265 ;
    END
END OAI222_X4_18_SVT_WB

MACRO OAI222_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI222_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.915 1.770 5.460 2.180 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 2.320 4.185 2.660 ;
        RECT  3.860 1.620 4.185 2.660 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.160 1.770 2.660 2.200 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.640 3.450 1.980 ;
        RECT  2.940 1.640 3.220 2.150 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.640 1.720 2.310 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.735 1.020 2.205 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.407  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.690 2.985 5.420 3.325 ;
        RECT  4.415 2.515 5.420 3.325 ;
        RECT  4.415 1.100 4.685 3.325 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  3.600 3.555 3.940 4.100 ;
        RECT  0.470 2.435 0.810 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  0.180 -0.180 0.520 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.685 1.240 1.410 ;
        RECT  0.900 1.070 3.260 1.410 ;
        RECT  2.200 0.565 5.420 0.840 ;
        RECT  3.640 0.565 3.980 1.375 ;
        RECT  5.080 0.565 5.420 1.385 ;
    END
END OAI222_X2_18_SVT_WB

MACRO OAI222_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI222_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.525 1.690 4.900 2.500 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.210 2.380 3.830 2.710 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.035 1.660 2.695 2.430 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.925 1.620 3.515 2.150 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.550 1.780 2.310 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.910 0.755 2.720 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.870  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.680 2.940 4.730 3.280 ;
        RECT  4.060 0.995 4.295 3.280 ;
        RECT  3.960 0.995 4.295 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.160 3.510 3.500 4.100 ;
        RECT  0.490 3.045 0.830 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  0.340 -0.180 1.720 0.465 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.790 0.980 2.980 1.320 ;
    END
END OAI222_X1_18_SVT_WB

MACRO OAI222_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI222_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.450 1.585 4.900 2.395 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.205 2.380 3.640 2.815 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.660 2.280 2.150 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.770 1.695 3.270 2.100 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.170  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.365 1.660 2.815 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.170  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 2.030 0.980 2.840 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 3.045 4.650 3.340 ;
        RECT  3.880 2.940 4.650 3.340 ;
        RECT  3.880 1.065 4.220 3.340 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.080 3.570 3.420 4.100 ;
        RECT  0.270 3.070 0.610 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.210 -0.180 1.550 0.560 ;
        RECT  0.180 -0.180 0.980 0.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.065 2.900 1.405 ;
    END
END OAI222_X0_18_SVT_WB

MACRO OAI221_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI221_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.385 1.445 7.695 2.065 ;
        RECT  5.175 1.445 7.695 1.675 ;
        RECT  5.175 1.445 6.060 2.185 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.290 1.905 6.670 2.720 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.770 2.980 2.060 ;
        RECT  2.380 1.410 2.685 2.060 ;
        RECT  0.435 1.410 2.685 1.640 ;
        RECT  0.435 1.410 1.050 2.150 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.660 2.250 2.225 2.660 ;
        RECT  1.660 1.915 2.050 2.660 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.345 1.805 4.800 2.185 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.925 0.985 8.260 2.830 ;
        RECT  0.175 3.030 8.010 3.305 ;
        RECT  7.585 2.480 8.010 3.305 ;
        RECT  5.195 0.985 8.260 1.215 ;
        RECT  0.175 3.015 5.750 3.305 ;
        RECT  4.855 2.905 5.750 3.305 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  6.355 3.560 6.705 4.100 ;
        RECT  4.155 3.560 4.515 4.100 ;
        RECT  1.525 3.570 1.865 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  2.840 -0.180 3.185 0.355 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.715 0.470 1.095 1.165 ;
        RECT  2.050 0.470 2.465 1.165 ;
        RECT  0.715 0.830 2.465 1.165 ;
        RECT  0.715 0.895 3.240 1.165 ;
        RECT  3.000 0.895 3.240 1.520 ;
        RECT  4.320 1.095 4.615 1.520 ;
        RECT  3.000 1.250 4.615 1.520 ;
        RECT  3.735 0.470 8.225 0.755 ;
        RECT  3.735 0.470 4.010 1.020 ;
        RECT  3.550 0.765 4.010 1.020 ;
    END
END OAI221_X4_18_SVT_WB

MACRO OAI221_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI221_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.210 4.340 1.590 ;
        RECT  3.750 1.210 4.090 2.060 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.740 3.060 2.080 ;
        RECT  2.620 1.260 2.850 2.080 ;
        RECT  2.330 1.260 2.850 1.600 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.690 1.720 2.150 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.355 1.135 2.660 ;
        RECT  0.650 1.860 1.000 2.660 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.380 2.390 2.660 ;
        RECT  2.050 1.860 2.390 2.660 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.740  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.620 3.045 3.970 3.280 ;
        RECT  3.290 2.940 3.970 3.280 ;
        RECT  3.290 1.100 3.520 3.280 ;
        RECT  3.080 1.100 3.520 1.440 ;
        RECT  1.620 3.045 1.960 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  2.380 3.515 2.720 4.100 ;
        RECT  0.470 3.110 0.810 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  0.900 -0.180 1.240 0.770 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.160 0.525 0.520 1.285 ;
        RECT  1.620 0.525 1.980 1.285 ;
        RECT  0.160 1.000 1.980 1.285 ;
        RECT  2.340 0.480 4.120 0.820 ;
    END
END OAI221_X2_18_SVT_WB

MACRO OAI221_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI221_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.060 3.805 2.060 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.770 2.725 2.330 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.665 1.390 2.150 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.565 2.380 1.190 2.730 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.685 2.190 2.115 2.710 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.870  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.520 2.940 3.730 3.245 ;
        RECT  2.955 2.925 3.730 3.245 ;
        RECT  2.955 1.005 3.185 3.245 ;
        RECT  2.720 1.005 3.185 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.350 2.990 0.690 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.800 -0.180 1.140 1.305 ;
        END
    END VSS
END OAI221_X1_18_SVT_WB

MACRO OAI221_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI221_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.400 1.750 3.790 2.560 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.335 1.620 2.710 2.160 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.950 1.540 2.710 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.345 1.770 0.670 2.760 ;
        RECT  0.115 1.770 0.670 2.395 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.370 2.190 2.710 ;
        RECT  1.770 2.180 2.105 2.710 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.370 2.940 3.580 3.280 ;
        RECT  2.940 1.100 3.170 3.280 ;
        RECT  2.810 1.100 3.170 1.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.220 2.995 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.890 -0.180 1.230 1.440 ;
        END
    END VSS
END OAI221_X0_18_SVT_WB

MACRO OAI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.523  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.970 1.370 4.390 2.130 ;
        RECT  1.740 1.370 4.390 1.600 ;
        RECT  1.740 1.370 2.080 2.005 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.523  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.620 1.720 5.605 2.060 ;
        RECT  1.235 2.690 4.935 2.920 ;
        RECT  4.620 1.720 4.935 2.920 ;
        RECT  2.580 1.905 2.920 2.920 ;
        RECT  1.235 1.875 1.510 2.920 ;
        RECT  0.575 1.875 1.510 2.300 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.955 1.695 7.175 2.230 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.618  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.620 2.695 7.960 3.450 ;
        RECT  6.180 1.080 7.960 1.385 ;
        RECT  7.405 1.080 7.765 2.925 ;
        RECT  5.570 2.695 7.960 2.925 ;
        RECT  1.500 3.150 5.800 3.380 ;
        RECT  5.570 2.695 5.800 3.380 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.340 2.640 8.680 4.100 ;
        RECT  6.900 3.165 7.240 4.100 ;
        RECT  0.350 2.530 0.690 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  3.570 -0.180 3.925 0.390 ;
        RECT  0.740 -0.180 1.080 0.360 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  5.460 0.510 8.680 0.850 ;
        RECT  5.460 0.510 5.785 1.130 ;
        RECT  0.180 0.890 5.785 1.130 ;
        RECT  8.340 0.510 8.680 1.320 ;
    END
END OAI21_X8_18_SVT_WB

MACRO OAI21_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.455 4.390 2.150 ;
        RECT  1.390 1.455 4.390 1.685 ;
        RECT  1.390 1.455 2.200 1.905 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.960 2.135 3.370 2.365 ;
        RECT  2.560 1.915 3.370 2.365 ;
        RECT  0.650 1.820 1.160 2.265 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.620 1.620 5.105 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.268  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.335 1.520 7.080 1.750 ;
        RECT  6.740 0.590 7.080 1.750 ;
        RECT  5.945 2.595 6.350 3.385 ;
        RECT  5.720 1.520 6.030 2.825 ;
        RECT  1.620 2.595 6.350 2.825 ;
        RECT  5.335 1.520 6.030 1.755 ;
        RECT  5.335 1.005 5.640 1.755 ;
        RECT  4.290 2.595 4.630 3.405 ;
        RECT  1.620 2.595 1.960 3.350 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.740 2.630 7.100 4.100 ;
        RECT  5.280 3.055 5.620 4.100 ;
        RECT  2.920 3.055 3.260 4.100 ;
        RECT  0.460 2.565 0.800 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  3.820 -0.180 4.160 0.405 ;
        RECT  2.340 -0.180 2.680 0.765 ;
        RECT  0.900 -0.180 1.240 0.765 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  4.580 0.535 6.360 0.775 ;
        RECT  3.060 0.525 3.400 1.225 ;
        RECT  0.180 0.525 0.520 1.225 ;
        RECT  1.620 0.525 1.960 1.225 ;
        RECT  3.060 0.885 4.920 1.225 ;
        RECT  0.180 0.995 4.920 1.225 ;
        RECT  6.020 0.535 6.360 1.290 ;
        RECT  4.580 0.535 4.920 1.315 ;
    END
END OAI21_X6_18_SVT_WB

MACRO OAI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.915 2.190 2.185 ;
        RECT  1.260 1.915 1.655 2.710 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.640 2.920 1.970 ;
        RECT  0.650 1.455 2.905 1.685 ;
        RECT  0.650 1.455 1.030 2.100 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.445 1.760 3.825 2.315 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.809  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.780 2.575 4.285 3.385 ;
        RECT  4.055 1.040 4.285 3.385 ;
        RECT  3.780 1.040 4.285 1.380 ;
        RECT  1.620 2.940 4.285 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.515 2.615 4.840 4.100 ;
        RECT  3.020 3.515 3.360 4.100 ;
        RECT  0.460 2.545 0.800 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  2.340 -0.180 2.680 0.765 ;
        RECT  0.900 -0.180 1.240 0.765 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.060 0.470 4.840 0.810 ;
        RECT  0.180 0.525 0.520 1.225 ;
        RECT  1.620 0.525 1.960 1.225 ;
        RECT  3.060 0.470 3.400 1.225 ;
        RECT  0.180 0.995 3.400 1.225 ;
        RECT  4.515 0.470 4.840 1.280 ;
    END
END OAI21_X4_18_SVT_WB

MACRO OAI21_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.596  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.410 2.065 2.220 2.765 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.596  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.550 1.595 2.890 1.935 ;
        RECT  0.650 1.595 2.890 1.835 ;
        RECT  0.650 1.595 1.030 2.100 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.596  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.095 1.770 4.900 2.165 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.361  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.625 3.010 4.140 3.340 ;
        RECT  3.405 2.780 4.140 3.340 ;
        RECT  3.635 1.005 4.140 1.345 ;
        RECT  3.635 1.005 3.865 3.340 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.520 3.030 4.860 4.100 ;
        RECT  2.830 3.570 3.170 4.100 ;
        RECT  0.490 2.585 0.830 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  2.360 -0.180 2.700 0.905 ;
        RECT  0.920 -0.180 1.260 0.905 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.080 0.410 4.860 0.750 ;
        RECT  4.520 0.410 4.860 0.975 ;
        RECT  0.200 0.635 0.540 1.365 ;
        RECT  1.640 1.005 1.980 1.365 ;
        RECT  3.080 0.410 3.405 1.365 ;
        RECT  0.200 1.135 3.405 1.365 ;
    END
END OAI21_X3_18_SVT_WB

MACRO OAI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.620 1.665 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.640 1.645 0.980 2.250 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.360 1.915 2.750 2.710 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.125  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.900 1.455 2.750 1.685 ;
        RECT  2.370 0.610 2.750 1.685 ;
        RECT  1.900 1.455 2.130 2.815 ;
        RECT  1.620 2.475 1.960 3.175 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.365 2.990 2.720 4.100 ;
        RECT  0.470 2.640 0.810 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.900 -0.180 1.240 0.765 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.525 0.520 1.225 ;
        RECT  1.620 0.525 1.960 1.225 ;
        RECT  0.180 0.995 1.960 1.225 ;
    END
END OAI21_X2_18_SVT_WB

MACRO OAI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 2.235 1.590 2.700 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.220 0.735 2.750 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.590 2.105 2.235 ;
        RECT  1.490 1.590 2.105 1.995 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.597  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.830 2.465 2.660 2.695 ;
        RECT  2.335 1.000 2.660 2.695 ;
        RECT  1.560 2.970 2.060 3.200 ;
        RECT  1.830 2.465 2.060 3.200 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.290 2.925 2.625 4.100 ;
        RECT  0.220 2.980 0.565 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.735 -0.180 1.090 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.055 1.840 1.285 ;
    END
END OAI21_X1_18_SVT_WB

MACRO OAI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.645 1.540 2.410 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.995 0.730 2.805 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.620 2.200 2.410 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.640 2.660 2.870 ;
        RECT  2.430 0.560 2.660 2.870 ;
        RECT  2.280 0.560 2.660 1.390 ;
        RECT  1.260 2.640 1.720 3.325 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.140 3.100 2.480 4.100 ;
        RECT  0.180 3.035 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.330 -0.180 1.140 0.650 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.045 1.900 1.390 ;
    END
END OAI21_X0_18_SVT_WB

MACRO OAI21P2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21P2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.161  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.010 1.390 3.830 2.110 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.110  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.435 2.195 2.100 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.110  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.510 1.500 5.225 2.140 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.991  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.220 2.380 7.170 2.720 ;
        RECT  6.825 0.845 7.170 2.720 ;
        RECT  5.455 1.365 7.170 1.595 ;
        RECT  5.455 0.870 5.725 1.595 ;
        RECT  5.370 0.870 5.725 1.160 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  6.825 2.950 7.165 4.100 ;
        RECT  5.385 3.110 5.725 4.100 ;
        RECT  1.625 3.110 1.965 4.100 ;
        RECT  0.185 3.110 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  2.465 -0.180 2.805 0.405 ;
        RECT  0.945 -0.180 1.285 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.905 2.640 2.845 2.880 ;
        RECT  2.505 2.640 2.845 3.450 ;
        RECT  0.905 2.640 1.245 3.450 ;
        RECT  2.505 3.110 4.285 3.450 ;
        RECT  4.665 0.410 6.445 0.640 ;
        RECT  4.665 0.410 5.005 0.990 ;
        RECT  0.185 0.650 5.005 0.990 ;
        RECT  6.105 0.410 6.445 0.990 ;
    END
END OAI21P2_X6_18_SVT_WB

MACRO OAI21P2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21P2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.635 1.540 2.275 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.720 2.160 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.670 2.140 2.320 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.858  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.370 3.060 2.660 3.400 ;
        RECT  2.370 1.100 2.660 3.400 ;
        RECT  2.280 1.100 2.660 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.165 2.990 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.860 -0.180 1.200 1.405 ;
        END
    END VSS
END OAI21P2_X1_18_SVT_WB

MACRO OAI21P2_X14_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21P2_X14_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.652  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.275 1.390 10.305 2.110 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.609  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.920 1.435 5.185 2.100 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.609  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.535 1.585 13.540 2.140 ;
        RECT  10.535 1.500 11.250 2.140 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.703  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.210 2.380 16.075 2.720 ;
        RECT  15.730 0.845 16.075 2.720 ;
        RECT  11.480 1.125 16.075 1.355 ;
        RECT  14.975 2.380 15.400 3.315 ;
        RECT  14.275 0.870 14.630 1.355 ;
        RECT  13.525 2.380 13.955 3.335 ;
        RECT  12.815 0.870 13.225 1.355 ;
        RECT  12.080 2.380 12.520 3.410 ;
        RECT  11.350 0.870 11.775 1.170 ;
        RECT  10.625 2.380 11.085 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  15.720 3.125 16.060 4.100 ;
        RECT  14.280 3.125 14.620 4.100 ;
        RECT  12.840 3.125 13.180 4.100 ;
        RECT  11.400 3.110 11.740 4.100 ;
        RECT  4.760 3.110 5.100 4.100 ;
        RECT  3.240 3.110 3.580 4.100 ;
        RECT  1.800 3.110 2.140 4.100 ;
        RECT  0.280 3.110 0.620 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  9.920 -0.180 10.260 0.350 ;
        RECT  6.960 -0.180 7.300 0.350 ;
        RECT  4.000 -0.180 4.340 0.350 ;
        RECT  1.040 -0.180 1.380 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.080 2.640 5.820 2.880 ;
        RECT  5.480 2.640 5.820 3.450 ;
        RECT  1.080 2.640 1.420 3.450 ;
        RECT  2.520 2.640 2.860 3.450 ;
        RECT  4.040 2.640 4.380 3.450 ;
        RECT  5.480 3.110 10.300 3.450 ;
        RECT  10.680 0.410 15.340 0.640 ;
        RECT  0.280 0.580 11.020 0.890 ;
        RECT  12.120 0.410 12.460 0.895 ;
        RECT  13.560 0.410 13.900 0.895 ;
        RECT  15.000 0.410 15.340 0.895 ;
    END
END OAI21P2_X14_18_SVT_WB

MACRO OAI21P2_X10_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21P2_X10_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.908  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.360 1.600 7.245 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.861  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.765 1.600 3.345 2.105 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.861  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.075 1.600 10.655 2.100 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.580 2.330 11.540 2.670 ;
        RECT  11.200 0.840 11.540 2.670 ;
        RECT  8.240 1.135 11.540 1.365 ;
        RECT  10.480 2.330 10.820 3.135 ;
        RECT  4.580 2.330 10.820 2.675 ;
        RECT  9.680 0.895 10.020 1.365 ;
        RECT  8.960 2.330 9.300 3.135 ;
        RECT  8.240 0.895 8.580 1.365 ;
        RECT  7.520 2.330 7.860 3.135 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  11.200 3.015 11.600 4.100 ;
        RECT  9.720 2.905 10.060 4.100 ;
        RECT  8.240 3.125 8.580 4.100 ;
        RECT  3.060 3.110 3.400 4.100 ;
        RECT  1.620 3.110 1.960 4.100 ;
        RECT  0.180 2.595 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  6.760 -0.180 7.100 0.410 ;
        RECT  3.820 -0.180 4.160 0.410 ;
        RECT  0.940 -0.180 1.280 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.640 4.200 2.880 ;
        RECT  3.860 2.640 4.200 3.450 ;
        RECT  0.900 2.640 1.240 3.395 ;
        RECT  2.340 2.640 2.680 3.395 ;
        RECT  3.860 3.110 7.080 3.450 ;
        RECT  7.520 0.435 10.740 0.665 ;
        RECT  8.960 0.435 9.300 0.905 ;
        RECT  10.400 0.435 10.740 0.905 ;
        RECT  7.520 0.435 7.860 1.030 ;
        RECT  0.180 0.690 7.860 1.030 ;
    END
END OAI21P2_X10_18_SVT_WB

MACRO OAI21P2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI21P2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.200 2.340 1.715 2.680 ;
        RECT  1.340 1.935 1.715 2.680 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.765 1.090 2.120 ;
        RECT  0.520 1.765 0.970 2.600 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.210 2.225 1.710 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.580 2.910 2.685 3.450 ;
        RECT  2.455 0.680 2.685 3.450 ;
        RECT  2.165 2.665 2.685 3.450 ;
        RECT  2.180 0.680 2.685 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.420 3.165 0.760 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.860 -0.180 1.200 1.440 ;
        END
    END VSS
END OAI21P2_X0_18_SVT_WB

MACRO OAI211_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI211_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.015 1.745 1.590 2.270 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.336  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.695 0.785 2.255 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.260 2.150 1.540 ;
        RECT  1.820 1.260 2.050 2.060 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.685 2.765 2.300 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.745 2.545 7.085 3.385 ;
        RECT  5.425 1.055 7.085 1.350 ;
        RECT  6.745 0.535 7.085 1.350 ;
        RECT  5.425 2.545 7.085 2.940 ;
        RECT  6.220 1.055 6.595 2.940 ;
        RECT  5.425 0.590 5.775 1.350 ;
        RECT  5.425 2.545 5.765 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  4.660 3.570 5.000 4.100 ;
        RECT  0.235 2.640 0.465 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  4.660 -0.180 5.000 0.350 ;
        RECT  0.820 -0.180 1.050 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.800 1.865 1.030 ;
        RECT  0.180 0.800 0.465 1.145 ;
        RECT  2.855 0.495 3.225 1.305 ;
        RECT  2.995 1.750 4.220 2.175 ;
        RECT  1.385 2.640 3.225 3.220 ;
        RECT  1.385 2.640 1.615 3.450 ;
        RECT  2.995 0.495 3.225 3.450 ;
        RECT  2.650 2.640 3.225 3.450 ;
        RECT  4.100 0.905 4.785 1.160 ;
        RECT  4.450 0.905 4.785 2.670 ;
        RECT  4.450 1.620 5.965 1.960 ;
        RECT  4.450 1.620 4.790 2.670 ;
        RECT  4.100 2.405 4.790 2.670 ;
    END
END OAI211_X8_18_SVT_WB

MACRO OAI211_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI211_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.815 1.585 2.710 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.410 1.260 2.695 2.060 ;
        RECT  0.275 1.260 2.695 1.540 ;
        RECT  0.275 1.260 0.595 2.080 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.490 2.460 5.560 2.690 ;
        RECT  5.230 1.260 5.560 2.690 ;
        RECT  5.115 1.260 5.560 1.625 ;
        RECT  3.490 1.555 3.720 2.690 ;
        RECT  3.385 1.555 3.720 2.060 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.865 4.830 2.180 ;
        RECT  4.060 1.670 4.360 2.180 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.518  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.010 3.045 5.350 3.385 ;
        RECT  1.500 3.045 5.350 3.285 ;
        RECT  2.925 1.095 4.595 1.325 ;
        RECT  3.490 3.045 3.830 3.385 ;
        RECT  1.500 2.940 3.155 3.285 ;
        RECT  2.925 1.095 3.155 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  2.730 3.515 3.070 4.100 ;
        RECT  0.180 2.640 0.500 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  2.260 -0.180 2.600 0.360 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.535 0.520 0.865 ;
        RECT  3.020 0.525 5.780 0.865 ;
        RECT  0.180 0.590 5.780 0.865 ;
    END
END OAI211_X4_18_SVT_WB

MACRO OAI211_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI211_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.015 1.745 1.590 2.270 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.336  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.695 0.785 2.255 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.260 2.150 1.540 ;
        RECT  1.820 1.260 2.050 2.060 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.685 2.765 2.300 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.677  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.650 2.640 3.225 3.450 ;
        RECT  2.995 0.495 3.225 3.450 ;
        RECT  2.855 0.495 3.225 1.305 ;
        RECT  1.385 2.640 3.225 3.220 ;
        RECT  1.385 2.640 1.615 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.235 2.640 0.465 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.820 -0.180 1.050 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.800 1.865 1.030 ;
        RECT  0.180 0.800 0.465 1.145 ;
    END
END OAI211_X2_18_SVT_WB

MACRO OAI211_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI211_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.955 1.540 2.765 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.490 2.300 0.980 2.710 ;
        RECT  0.490 1.540 0.830 2.710 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.190 2.255 1.615 ;
        RECT  1.820 1.190 2.150 2.470 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.955 2.785 2.765 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.839  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.740 2.995 3.245 3.335 ;
        RECT  3.015 0.645 3.245 3.335 ;
        RECT  2.740 0.645 3.245 1.030 ;
        RECT  1.400 2.995 3.245 3.320 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.250 3.035 0.590 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.415 -0.180 1.115 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.590 0.540 1.930 0.960 ;
        RECT  0.250 0.730 1.930 0.960 ;
        RECT  0.250 0.730 0.590 1.305 ;
    END
END OAI211_X1_18_SVT_WB

MACRO OAI211_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI211_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.580 1.550 2.805 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.635 0.980 2.150 ;
        RECT  0.490 1.635 0.830 2.805 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.815 1.160 2.275 1.600 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.350 2.050 2.690 2.810 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.400 3.040 3.220 3.380 ;
        RECT  2.920 0.590 3.220 3.380 ;
        RECT  2.840 0.590 3.220 0.930 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.250 3.095 0.590 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.515 -0.180 1.215 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.690 0.590 2.030 0.930 ;
        RECT  0.240 0.700 2.030 0.930 ;
        RECT  0.240 0.700 0.580 1.350 ;
    END
END OAI211_X0_18_SVT_WB

MACRO OAI12_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 1.455 5.015 2.110 ;
        RECT  2.125 1.455 5.015 1.685 ;
        RECT  2.125 1.455 2.460 1.980 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.920 2.345 6.145 2.670 ;
        RECT  5.800 1.670 6.145 2.670 ;
        RECT  0.920 2.330 3.675 2.670 ;
        RECT  3.335 1.915 3.675 2.670 ;
        RECT  0.920 1.640 1.260 2.670 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.670 8.295 2.100 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.936  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.600 1.210 8.940 3.450 ;
        RECT  7.030 2.650 8.940 2.880 ;
        RECT  8.595 1.210 8.940 2.880 ;
        RECT  5.560 1.210 8.940 1.440 ;
        RECT  7.065 2.650 7.520 3.440 ;
        RECT  1.880 2.940 7.520 3.280 ;
        RECT  7.030 2.650 7.520 3.280 ;
        RECT  1.160 0.995 5.920 1.225 ;
        RECT  1.160 0.995 1.500 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  9.320 2.640 9.660 4.100 ;
        RECT  7.880 3.110 8.220 4.100 ;
        RECT  6.115 3.515 6.455 4.100 ;
        RECT  3.360 3.515 3.700 4.100 ;
        RECT  0.440 3.110 0.730 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  8.560 -0.180 8.900 0.405 ;
        RECT  7.040 -0.180 7.380 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.440 0.470 6.620 0.765 ;
        RECT  6.280 0.645 9.660 0.975 ;
        RECT  0.440 0.470 0.780 1.280 ;
    END
END OAI12_X8_18_SVT_WB

MACRO OAI12_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.810 4.120 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.760 1.805 2.100 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.000 1.680 6.300 2.100 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.656  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.960 2.380 6.300 3.230 ;
        RECT  3.080 2.380 6.300 2.720 ;
        RECT  4.350 1.105 4.690 2.720 ;
        RECT  0.920 1.105 4.690 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.760 2.450 7.100 4.100 ;
        RECT  5.240 3.110 5.580 4.100 ;
        RECT  1.640 3.110 1.980 4.100 ;
        RECT  0.200 2.600 0.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.760 -0.180 7.100 1.345 ;
        RECT  5.280 -0.180 5.620 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.920 2.380 2.700 2.720 ;
        RECT  2.360 2.380 2.700 3.235 ;
        RECT  0.920 2.380 1.260 3.190 ;
        RECT  2.360 2.950 4.140 3.235 ;
        RECT  0.200 0.535 4.860 0.875 ;
        RECT  6.040 0.535 6.380 0.875 ;
        RECT  0.200 0.635 6.380 0.875 ;
        RECT  0.200 0.535 0.540 1.440 ;
    END
END OAI12_X6_18_SVT_WB

MACRO OAI12_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.640 3.470 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.170 2.330 4.360 2.670 ;
        RECT  4.020 1.620 4.360 2.670 ;
        RECT  2.170 1.640 2.510 2.670 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.605 1.620 1.030 2.100 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.920 2.945 4.925 3.285 ;
        RECT  4.590 1.040 4.925 3.285 ;
        RECT  2.360 1.040 4.925 1.380 ;
        RECT  0.920 2.475 1.260 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.270 3.515 4.610 4.100 ;
        RECT  1.890 3.515 2.230 4.100 ;
        RECT  0.200 2.475 0.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  0.920 -0.180 1.260 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.640 0.470 4.860 0.810 ;
        RECT  0.200 0.470 0.540 1.280 ;
        RECT  1.640 0.470 1.980 1.280 ;
        RECT  0.200 1.040 1.980 1.280 ;
    END
END OAI12_X4_18_SVT_WB

MACRO OAI12_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.596  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.820 1.665 3.240 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.596  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.150 2.380 4.340 2.705 ;
        RECT  4.000 1.560 4.340 2.705 ;
        RECT  2.150 2.005 2.490 2.705 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.596  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 1.690 1.115 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.787  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 1.100 4.120 1.330 ;
        RECT  3.780 0.990 4.120 1.330 ;
        RECT  0.900 2.940 3.400 3.280 ;
        RECT  2.340 0.990 2.680 1.330 ;
        RECT  1.580 1.545 2.590 1.775 ;
        RECT  2.340 0.990 2.590 1.775 ;
        RECT  1.580 1.545 1.920 3.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.210 2.940 4.550 4.100 ;
        RECT  1.870 3.515 2.210 4.100 ;
        RECT  0.180 2.940 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  0.900 -0.180 1.240 0.855 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.620 0.530 4.840 0.760 ;
        RECT  3.060 0.530 3.400 0.870 ;
        RECT  4.500 0.530 4.840 0.925 ;
        RECT  0.180 0.585 0.520 1.315 ;
        RECT  1.620 0.530 1.960 1.315 ;
        RECT  0.180 1.085 1.960 1.315 ;
    END
END OAI12_X3_18_SVT_WB

MACRO OAI12_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.545 1.655 2.100 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.670 0.505 2.260 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.640 2.730 2.145 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 2.380 2.190 3.310 ;
        RECT  1.085 2.380 2.190 2.840 ;
        RECT  1.085 1.085 1.470 1.425 ;
        RECT  1.085 1.085 1.315 2.840 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.570 2.500 2.910 4.100 ;
        RECT  0.410 2.490 0.750 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.570 -0.180 2.910 1.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.410 0.615 2.190 0.855 ;
        RECT  1.850 0.615 2.190 1.425 ;
        RECT  0.410 0.615 0.750 1.440 ;
    END
END OAI12_X2_18_SVT_WB

MACRO OAI12_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.595 1.590 2.250 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.570 2.345 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.725 2.295 2.155 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.800 2.520 1.805 2.920 ;
        RECT  0.800 0.970 1.030 2.920 ;
        RECT  0.500 1.250 1.030 1.540 ;
        RECT  0.710 0.970 1.030 1.540 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.185 2.535 2.525 4.100 ;
        RECT  0.275 2.990 0.570 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.185 -0.180 2.525 1.415 ;
        END
    END VSS
END OAI12_X1_18_SVT_WB

MACRO OAI12_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.600 2.290 2.150 2.660 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.525 0.655 2.415 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.770 2.915 2.110 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 2.890 2.160 3.230 ;
        RECT  1.100 1.100 1.440 1.900 ;
        RECT  1.100 1.100 1.370 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.540 2.890 2.880 4.100 ;
        RECT  0.380 2.890 0.720 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.540 -0.180 2.880 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.340 0.630 2.160 0.870 ;
        RECT  0.340 0.630 0.680 0.970 ;
        RECT  1.820 0.630 2.160 1.440 ;
    END
END OAI12_X0_18_SVT_WB

MACRO OAI12P2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12P2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.156  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.740 1.575 3.555 2.120 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.106  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.980 1.560 1.950 2.125 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.106  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.060 1.575 6.600 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.406  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.965 2.380 6.360 3.450 ;
        RECT  3.860 2.380 6.360 2.610 ;
        RECT  4.580 2.380 4.920 3.385 ;
        RECT  3.140 2.570 4.920 2.910 ;
        RECT  3.860 0.870 4.200 2.910 ;
        RECT  0.900 1.100 4.200 1.330 ;
        RECT  2.420 0.870 2.760 1.330 ;
        RECT  0.900 0.870 1.240 1.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.740 2.600 7.080 4.100 ;
        RECT  5.300 3.095 5.640 4.100 ;
        RECT  1.660 3.515 2.000 4.100 ;
        RECT  0.180 2.575 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.740 -0.180 7.080 1.095 ;
        RECT  5.300 -0.180 5.640 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.575 2.760 2.805 ;
        RECT  2.420 2.575 2.760 3.425 ;
        RECT  0.900 2.575 1.240 3.385 ;
        RECT  2.420 3.140 4.200 3.425 ;
        RECT  0.180 0.410 4.920 0.640 ;
        RECT  0.180 0.410 0.520 0.870 ;
        RECT  1.620 0.410 1.960 0.870 ;
        RECT  3.140 0.410 3.480 0.870 ;
        RECT  4.580 0.410 4.920 1.345 ;
        RECT  6.020 0.535 6.360 1.345 ;
        RECT  4.580 1.115 6.360 1.345 ;
    END
END OAI12P2_X6_18_SVT_WB

MACRO OAI12P2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12P2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.705 1.695 2.220 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.620 0.520 2.285 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.655 2.685 2.220 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.695 2.870 1.900 3.450 ;
        RECT  1.560 2.640 1.900 3.450 ;
        RECT  0.750 1.100 1.175 1.440 ;
        RECT  0.695 2.795 0.980 3.450 ;
        RECT  0.750 1.100 0.980 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.280 2.640 2.620 4.100 ;
        RECT  0.180 2.630 0.465 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.280 -0.180 2.620 1.425 ;
        END
    END VSS
END OAI12P2_X1_18_SVT_WB

MACRO OAI12P2_X14_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12P2_X14_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.640  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.980 1.560 8.800 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.598  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.560 4.305 2.150 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.598  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.090 1.475 14.880 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.868  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.000 2.415 14.980 2.720 ;
        RECT  11.760 2.415 12.100 3.450 ;
        RECT  6.000 2.410 10.660 2.720 ;
        RECT  9.600 0.870 9.940 2.720 ;
        RECT  0.960 1.100 9.940 1.330 ;
        RECT  8.160 0.870 8.500 1.330 ;
        RECT  6.720 0.870 7.060 1.330 ;
        RECT  5.280 0.870 5.620 1.330 ;
        RECT  3.840 0.870 4.180 1.330 ;
        RECT  2.400 0.870 2.740 1.330 ;
        RECT  0.960 0.870 1.300 1.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  15.360 2.600 15.700 4.100 ;
        RECT  13.920 3.110 14.260 4.100 ;
        RECT  12.480 3.110 12.820 4.100 ;
        RECT  11.040 3.110 11.380 4.100 ;
        RECT  4.560 3.110 4.900 4.100 ;
        RECT  3.120 3.110 3.460 4.100 ;
        RECT  1.680 3.110 2.020 4.100 ;
        RECT  0.240 2.380 0.580 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  15.600 -0.180 15.940 0.980 ;
        RECT  14.120 -0.180 14.460 0.420 ;
        RECT  12.600 -0.180 12.940 0.420 ;
        RECT  11.080 -0.180 11.420 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.960 2.380 5.620 2.620 ;
        RECT  5.280 2.380 5.620 3.450 ;
        RECT  0.960 2.380 1.300 3.450 ;
        RECT  2.400 2.380 2.740 3.450 ;
        RECT  3.840 2.380 4.180 3.450 ;
        RECT  5.280 3.110 9.940 3.450 ;
        RECT  0.240 0.410 10.660 0.640 ;
        RECT  10.320 0.410 10.660 1.200 ;
        RECT  1.680 0.410 2.020 0.870 ;
        RECT  3.120 0.410 3.460 0.870 ;
        RECT  4.560 0.410 4.900 0.870 ;
        RECT  6.000 0.410 6.340 0.870 ;
        RECT  7.440 0.410 7.780 0.870 ;
        RECT  8.880 0.410 9.220 0.870 ;
        RECT  0.240 0.410 0.580 0.915 ;
        RECT  10.320 0.860 15.220 1.200 ;
    END
END OAI12P2_X14_18_SVT_WB

MACRO OAI12P2_X10_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12P2_X10_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.895  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.000 1.615 6.220 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.850  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 1.615 3.350 2.100 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.850  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.985 1.615 10.220 2.100 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.500 2.595 10.600 2.935 ;
        RECT  8.820 2.595 9.160 3.450 ;
        RECT  6.660 0.905 7.140 2.935 ;
        RECT  0.900 1.135 7.140 1.365 ;
        RECT  5.220 0.905 5.560 1.365 ;
        RECT  3.780 0.905 4.120 1.365 ;
        RECT  2.340 0.905 2.680 1.365 ;
        RECT  0.900 0.905 1.240 1.365 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  10.980 2.380 11.320 4.100 ;
        RECT  9.540 3.165 9.880 4.100 ;
        RECT  3.060 3.110 3.400 4.100 ;
        RECT  1.620 3.110 1.960 4.100 ;
        RECT  0.180 2.600 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  10.980 -0.180 11.320 0.975 ;
        RECT  9.540 -0.180 9.880 0.855 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.380 4.120 2.720 ;
        RECT  3.780 2.380 4.120 3.450 ;
        RECT  0.900 2.380 1.240 3.190 ;
        RECT  2.340 2.380 2.680 3.230 ;
        RECT  3.780 3.165 7.000 3.450 ;
        RECT  0.180 0.445 9.160 0.675 ;
        RECT  0.180 0.445 0.520 0.905 ;
        RECT  1.620 0.445 1.960 0.905 ;
        RECT  3.060 0.445 3.400 0.905 ;
        RECT  4.500 0.445 4.840 0.905 ;
        RECT  5.940 0.445 6.280 0.905 ;
        RECT  7.380 0.445 9.160 0.905 ;
        RECT  8.820 0.445 9.160 1.315 ;
        RECT  10.260 0.855 10.600 1.315 ;
        RECT  8.820 1.085 10.600 1.315 ;
    END
END OAI12P2_X10_18_SVT_WB

MACRO OAI12P2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OAI12P2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.770 1.670 2.280 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.210 0.470 2.015 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.060 1.720 2.660 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.680  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.510 1.900 2.850 ;
        RECT  0.700 1.100 1.180 1.440 ;
        RECT  0.700 1.100 1.020 2.850 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.280 2.905 2.620 4.100 ;
        RECT  0.370 3.480 0.710 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.280 -0.180 2.620 1.440 ;
        END
    END VSS
END OAI12P2_X0_18_SVT_WB

MACRO OA22_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA22_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.915 4.950 2.660 ;
        RECT  4.140 1.915 4.950 2.200 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.320 1.455 5.660 1.960 ;
        RECT  3.440 1.455 5.660 1.685 ;
        RECT  3.440 1.455 3.790 2.150 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.915 2.190 2.200 ;
        RECT  1.260 1.915 1.600 2.710 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.720 1.455 3.060 1.960 ;
        RECT  0.650 1.455 3.060 1.685 ;
        RECT  0.650 1.455 1.030 2.100 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.362  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.080 0.810 8.740 1.225 ;
        RECT  6.810 2.415 8.640 3.220 ;
        RECT  7.615 0.810 7.965 3.220 ;
        RECT  7.080 0.525 7.420 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  9.000 3.515 9.340 4.100 ;
        RECT  5.570 3.515 6.380 4.100 ;
        RECT  3.190 3.515 3.530 4.100 ;
        RECT  0.180 2.435 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  9.000 -0.180 9.340 0.405 ;
        RECT  0.900 -0.180 1.240 0.765 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.940 0.470 6.160 0.765 ;
        RECT  1.620 0.525 1.960 1.225 ;
        RECT  0.180 0.525 0.520 1.225 ;
        RECT  1.620 0.885 3.280 1.225 ;
        RECT  2.940 0.470 3.280 1.225 ;
        RECT  0.180 0.995 3.280 1.225 ;
        RECT  3.660 0.995 6.370 1.225 ;
        RECT  6.140 0.995 6.370 3.285 ;
        RECT  6.140 1.840 7.365 2.180 ;
        RECT  6.140 1.840 6.480 3.285 ;
        RECT  1.620 2.945 6.480 3.285 ;
    END
END OA22_X8_18_SVT_WB

MACRO OA22_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA22_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.710 1.720 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 1.620 1.000 2.215 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.255 1.620 2.710 2.100 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.760 3.500 2.150 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.395  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.375 2.875 4.900 3.385 ;
        RECT  4.375 0.535 4.700 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  5.130 2.575 5.420 4.100 ;
        RECT  3.390 3.100 3.775 4.100 ;
        RECT  0.180 2.435 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  5.080 -0.180 5.420 1.290 ;
        RECT  3.640 -0.180 3.980 0.875 ;
        RECT  2.160 -0.180 2.500 0.400 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.920 0.535 3.260 0.925 ;
        RECT  0.900 0.630 3.260 0.925 ;
        RECT  0.180 0.685 0.520 1.390 ;
        RECT  0.180 1.155 4.145 1.390 ;
        RECT  3.860 1.155 4.145 2.610 ;
        RECT  1.905 2.380 4.145 2.610 ;
        RECT  1.905 2.380 2.250 3.190 ;
    END
END OA22_X4_18_SVT_WB

MACRO OA22_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA22_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.184  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.760 1.455 3.100 ;
        RECT  1.170 2.240 1.455 3.100 ;
        RECT  0.700 2.760 1.040 3.330 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.179  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.500 2.070 0.840 2.530 ;
        RECT  0.140 2.070 0.840 2.300 ;
        RECT  0.140 1.645 0.480 2.300 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 1.770 2.660 2.580 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.770 3.225 2.580 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.995 2.480 4.340 3.435 ;
        RECT  4.060 0.595 4.340 3.435 ;
        RECT  3.995 0.595 4.340 1.425 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.200 3.515 3.540 4.100 ;
        RECT  0.185 2.760 0.470 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  2.040 -0.180 3.540 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.380 0.430 1.720 0.915 ;
        RECT  1.380 0.685 2.940 0.915 ;
        RECT  2.600 0.685 2.940 1.145 ;
        RECT  0.780 1.200 1.915 1.540 ;
        RECT  3.480 1.720 3.830 2.070 ;
        RECT  1.685 1.200 1.915 3.150 ;
        RECT  3.480 1.720 3.765 3.150 ;
        RECT  1.685 2.810 3.765 3.150 ;
    END
END OA22_X2_18_SVT_WB

MACRO OA22_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA22_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.245 2.305 1.665 2.850 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.152  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.075 0.785 2.480 ;
        RECT  0.140 1.760 0.465 2.480 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.260 2.340 1.615 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.770 1.635 3.220 2.390 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.000 0.805 4.340 3.115 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.195 3.495 3.555 4.100 ;
        RECT  0.300 2.805 0.710 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  2.060 -0.180 3.540 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.330 0.420 1.830 0.765 ;
        RECT  1.600 0.690 2.960 0.920 ;
        RECT  2.620 0.690 2.960 1.145 ;
        RECT  0.800 1.170 1.275 1.510 ;
        RECT  1.045 1.170 1.275 2.075 ;
        RECT  1.045 1.845 2.235 2.075 ;
        RECT  1.895 1.845 2.235 3.115 ;
        RECT  3.480 2.095 3.770 3.115 ;
        RECT  1.895 2.780 3.770 3.115 ;
    END
END OA22_X1_18_SVT_WB

MACRO OA22_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA22_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.125 1.710 2.725 2.125 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.635 3.780 2.390 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.715 2.355 2.355 2.755 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.690 1.680 2.110 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.480  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 0.470 1.090 0.980 ;
        RECT  0.115 2.795 0.600 3.080 ;
        RECT  0.115 0.470 0.345 3.080 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.415 2.990 3.740 4.100 ;
        RECT  0.820 3.565 1.160 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.450 -0.180 1.790 0.450 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.080 0.430 2.525 0.770 ;
        RECT  2.080 0.430 2.310 1.460 ;
        RECT  0.790 1.210 2.310 1.460 ;
        RECT  2.740 1.170 3.185 1.480 ;
        RECT  0.575 2.000 0.890 2.565 ;
        RECT  0.830 2.335 1.060 3.330 ;
        RECT  2.955 1.170 3.185 3.330 ;
        RECT  0.830 2.990 3.185 3.330 ;
    END
END OA22_X0_18_SVT_WB

MACRO OA21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.195  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.635 1.340 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.195  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.330 0.815 2.775 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.207  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.770 2.100 2.280 ;
        RECT  1.690 1.770 1.975 2.330 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.745 2.545 7.085 3.385 ;
        RECT  5.425 1.055 7.085 1.350 ;
        RECT  6.745 0.535 7.085 1.350 ;
        RECT  5.425 2.545 7.085 2.940 ;
        RECT  6.220 1.055 6.595 2.940 ;
        RECT  5.425 0.590 5.775 1.350 ;
        RECT  5.425 2.545 5.765 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  4.660 3.570 5.000 4.100 ;
        RECT  2.120 3.165 2.460 4.100 ;
        RECT  0.250 3.055 0.590 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  4.660 -0.180 5.000 0.350 ;
        RECT  2.120 -0.180 2.460 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.780 1.040 1.065 1.400 ;
        RECT  0.780 1.145 2.645 1.400 ;
        RECT  2.330 1.145 2.645 2.935 ;
        RECT  1.400 2.705 2.645 2.935 ;
        RECT  1.400 2.705 1.740 3.345 ;
        RECT  2.875 1.750 4.220 2.080 ;
        RECT  2.875 0.470 3.220 3.450 ;
        RECT  4.100 0.905 4.785 1.160 ;
        RECT  4.450 0.905 4.785 2.670 ;
        RECT  4.450 1.620 5.965 1.960 ;
        RECT  4.450 1.620 4.790 2.670 ;
        RECT  4.100 2.405 4.790 2.670 ;
    END
END OA21_X8_18_SVT_WB

MACRO OA21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.155 1.625 1.540 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.760 0.750 2.185 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.620 2.180 2.185 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.441  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.105 1.210 3.520 3.450 ;
        RECT  3.180 0.590 3.520 3.450 ;
        RECT  2.940 1.210 3.520 1.590 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.900 2.475 4.300 4.100 ;
        RECT  2.175 3.045 2.515 4.100 ;
        RECT  0.165 2.545 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.900 -0.180 4.300 1.345 ;
        RECT  2.420 -0.180 2.760 0.885 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 0.590 2.000 0.885 ;
        RECT  0.220 0.590 0.560 1.345 ;
        RECT  0.940 1.115 2.640 1.390 ;
        RECT  2.410 1.115 2.640 2.645 ;
        RECT  2.410 1.860 2.875 2.645 ;
        RECT  1.415 2.415 2.875 2.645 ;
        RECT  1.415 2.415 1.755 3.170 ;
    END
END OA21_X4_18_SVT_WB

MACRO OA21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.195  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.635 1.340 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.195  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.330 0.815 2.775 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.207  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.770 2.100 2.280 ;
        RECT  1.690 1.770 1.975 2.330 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.054  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.875 0.470 3.220 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.120 3.165 2.460 4.100 ;
        RECT  0.250 3.055 0.590 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.120 -0.180 2.460 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.780 1.040 1.065 1.400 ;
        RECT  0.780 1.145 2.645 1.400 ;
        RECT  2.330 1.145 2.645 2.935 ;
        RECT  1.400 2.705 2.645 2.935 ;
        RECT  1.400 2.705 1.740 3.345 ;
    END
END OA21_X2_18_SVT_WB

MACRO OA21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.255 1.610 1.540 2.150 ;
        RECT  0.925 1.610 1.540 1.950 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.435 2.380 1.030 2.720 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.385 2.100 2.725 ;
        RECT  1.770 1.965 2.100 2.725 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.880 0.580 3.220 2.825 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.335 3.425 3.035 4.100 ;
        RECT  0.325 3.010 0.710 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.120 -0.180 2.460 0.905 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.800 1.000 1.140 1.370 ;
        RECT  0.800 1.140 2.650 1.370 ;
        RECT  2.330 1.140 2.650 3.195 ;
        RECT  1.520 2.955 2.650 3.195 ;
        RECT  1.520 2.955 1.860 3.295 ;
    END
END OA21_X1_18_SVT_WB

MACRO OA21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN OA21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.980 1.645 1.740 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.560 0.760 2.865 ;
        RECT  0.140 2.105 0.600 2.865 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 2.380 2.150 2.865 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.855 0.540 3.220 3.435 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 3.095 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.120 -0.180 2.460 0.845 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.075 2.625 1.415 ;
        RECT  2.380 1.075 2.625 3.435 ;
        RECT  1.460 3.095 2.625 3.435 ;
    END
END OA21_X0_18_SVT_WB

MACRO NOR4_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR4_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.680 1.260 10.020 1.905 ;
        RECT  7.280 1.260 10.020 1.590 ;
        RECT  7.280 1.260 7.620 1.905 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.180 2.135 11.080 2.365 ;
        RECT  10.740 1.915 11.080 2.365 ;
        RECT  8.305 1.820 9.005 2.365 ;
        RECT  6.180 1.840 6.520 2.365 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.755 2.330 5.540 2.560 ;
        RECT  5.180 1.620 5.540 2.560 ;
        RECT  0.755 2.220 3.510 2.560 ;
        RECT  2.700 1.915 3.510 2.560 ;
        RECT  0.755 1.840 1.050 2.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.455 4.470 2.100 ;
        RECT  1.525 1.455 4.470 1.685 ;
        RECT  1.525 1.455 2.225 1.960 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.847  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.330 2.595 11.645 2.835 ;
        RECT  11.310 1.455 11.645 2.835 ;
        RECT  10.520 1.455 11.645 1.685 ;
        RECT  10.520 0.470 10.860 1.685 ;
        RECT  6.420 0.470 10.860 0.810 ;
        RECT  0.900 0.995 6.760 1.225 ;
        RECT  6.420 0.470 6.760 1.225 ;
        RECT  4.980 0.525 5.320 1.225 ;
        RECT  3.660 0.525 4.000 1.225 ;
        RECT  2.220 0.525 2.560 1.225 ;
        RECT  0.900 0.525 1.240 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  4.220 3.515 4.560 4.100 ;
        RECT  1.660 3.515 2.000 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  11.240 -0.180 11.580 1.225 ;
        RECT  5.700 -0.180 6.040 0.765 ;
        RECT  0.180 -0.180 0.520 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.295 2.395 0.525 3.285 ;
        RECT  0.295 3.000 5.065 3.285 ;
        RECT  4.725 3.065 11.300 3.350 ;
    END
END NOR4_X8_18_SVT_WB

MACRO NOR4_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR4_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.910 2.135 8.260 2.365 ;
        RECT  7.940 1.770 8.260 2.365 ;
        RECT  5.910 1.915 6.250 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.040 1.455 7.380 1.905 ;
        RECT  4.570 1.455 7.380 1.685 ;
        RECT  4.570 1.455 4.950 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.870 1.455 4.340 2.150 ;
        RECT  1.740 1.455 4.340 1.685 ;
        RECT  1.740 1.455 2.080 1.905 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 2.135 3.040 2.365 ;
        RECT  2.700 1.915 3.040 2.365 ;
        RECT  0.420 1.820 1.030 2.365 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.644  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.670 2.595 8.820 2.825 ;
        RECT  8.490 0.970 8.820 2.825 ;
        RECT  0.900 0.970 8.820 1.225 ;
        RECT  7.720 0.455 8.070 1.225 ;
        RECT  6.375 0.465 6.745 1.225 ;
        RECT  5.080 0.460 5.415 1.225 ;
        RECT  3.620 0.470 3.985 1.225 ;
        RECT  2.220 0.455 2.560 1.225 ;
        RECT  0.900 0.460 1.240 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  2.690 3.515 3.030 4.100 ;
        RECT  0.180 2.595 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.440 -0.180 8.780 0.740 ;
        RECT  4.350 -0.180 4.690 0.740 ;
        RECT  0.180 -0.180 0.520 1.305 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.500 2.595 3.580 2.935 ;
        RECT  3.240 2.595 3.580 3.395 ;
        RECT  3.240 3.055 7.160 3.395 ;
        RECT  1.500 2.595 1.860 3.465 ;
    END
END NOR4_X6_18_SVT_WB

MACRO NOR4_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR4_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.755 2.895 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.125 1.885 4.885 2.185 ;
        RECT  1.770 2.380 3.355 2.610 ;
        RECT  3.125 1.885 3.355 2.610 ;
        RECT  1.770 1.820 2.150 2.610 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.295 1.315 5.525 2.060 ;
        RECT  4.570 1.315 5.525 1.545 ;
        RECT  1.195 1.260 4.950 1.490 ;
        RECT  1.195 1.260 1.425 2.060 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.735 2.995 6.445 3.225 ;
        RECT  6.215 1.825 6.445 3.225 ;
        RECT  5.690 2.940 6.445 3.225 ;
        RECT  0.735 1.860 0.965 3.225 ;
        RECT  0.470 1.860 0.965 2.090 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.734  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.585 2.480 5.985 2.710 ;
        RECT  5.755 0.700 5.985 2.710 ;
        RECT  5.590 0.700 5.985 1.090 ;
        RECT  0.900 0.700 5.985 0.980 ;
        RECT  3.585 2.480 3.925 2.765 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  0.275 2.640 0.505 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  4.830 -0.180 5.060 0.405 ;
        RECT  3.180 -0.180 3.520 0.350 ;
        RECT  1.660 -0.180 2.000 0.350 ;
        RECT  0.235 -0.180 0.465 1.280 ;
        END
    END VSS
END NOR4_X4_18_SVT_WB

MACRO NOR4_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR4_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.510 2.765 2.330 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.620 2.150 2.170 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.575 1.540 2.395 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.705 0.760 2.220 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.697  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.720 2.560 3.225 3.260 ;
        RECT  2.995 0.470 3.225 3.260 ;
        RECT  2.205 0.470 3.225 1.280 ;
        RECT  0.900 0.470 3.225 0.755 ;
        RECT  0.900 0.470 1.240 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 2.450 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.180 -0.180 0.520 1.385 ;
        END
    END VSS
END NOR4_X2_18_SVT_WB

MACRO NOR4_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR4_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.705 2.720 2.515 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.955 2.150 2.765 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.485 1.540 2.150 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.190 2.380 1.030 2.785 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.843  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.670 2.890 3.220 3.285 ;
        RECT  2.950 0.860 3.220 3.285 ;
        RECT  0.900 0.860 3.220 1.200 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.420 3.100 0.760 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.825 -0.180 3.050 0.405 ;
        RECT  0.180 -0.180 0.520 1.200 ;
        END
    END VSS
END NOR4_X1_18_SVT_WB

MACRO NOR4_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR4_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.270 2.135 16.150 2.365 ;
        RECT  15.740 1.820 16.150 2.365 ;
        RECT  13.320 1.915 13.660 2.365 ;
        RECT  10.270 1.915 10.610 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.380 1.905 17.240 2.200 ;
        RECT  16.380 1.260 16.660 2.200 ;
        RECT  14.560 1.260 16.660 1.590 ;
        RECT  14.280 1.455 14.755 1.905 ;
        RECT  9.240 1.455 14.755 1.685 ;
        RECT  11.400 1.455 11.740 1.905 ;
        RECT  9.240 1.455 9.580 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.330 8.620 2.660 ;
        RECT  8.280 1.840 8.620 2.660 ;
        RECT  0.650 2.320 6.440 2.660 ;
        RECT  6.100 1.915 6.440 2.660 ;
        RECT  3.280 1.915 3.620 2.660 ;
        RECT  0.650 1.860 1.020 2.660 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.455 7.420 2.100 ;
        RECT  1.840 1.455 7.420 1.685 ;
        RECT  4.240 1.455 4.580 1.960 ;
        RECT  1.840 1.455 2.180 1.980 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 8.874  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.490 2.595 17.805 2.835 ;
        RECT  17.470 1.440 17.805 2.835 ;
        RECT  16.890 1.440 17.805 1.670 ;
        RECT  16.890 0.470 17.120 1.670 ;
        RECT  16.680 0.470 17.120 1.030 ;
        RECT  13.800 0.470 17.120 0.810 ;
        RECT  2.320 0.995 14.140 1.225 ;
        RECT  13.800 0.470 14.140 1.225 ;
        RECT  12.360 0.525 12.700 1.225 ;
        RECT  10.920 0.525 11.260 1.225 ;
        RECT  9.480 0.525 9.820 1.225 ;
        RECT  8.040 0.525 8.380 1.225 ;
        RECT  6.600 0.525 6.940 1.225 ;
        RECT  5.280 0.525 5.620 1.225 ;
        RECT  3.760 0.525 4.100 1.225 ;
        RECT  2.320 0.470 2.660 1.225 ;
        RECT  0.900 0.470 2.660 0.810 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  7.070 3.515 7.410 4.100 ;
        RECT  4.520 3.515 4.860 4.100 ;
        RECT  1.740 3.515 2.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  17.400 -0.180 17.740 1.210 ;
        RECT  13.080 -0.180 13.420 0.740 ;
        RECT  8.760 -0.180 9.100 0.765 ;
        RECT  4.520 -0.180 4.860 0.490 ;
        RECT  0.180 -0.180 0.520 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.460 2.990 8.155 3.285 ;
        RECT  7.815 3.065 17.460 3.350 ;
    END
END NOR4_X12_18_SVT_WB

MACRO NOR4_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR4_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.470 2.785 2.280 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 2.070 2.150 2.880 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.770 1.540 2.160 ;
        RECT  1.140 1.430 1.480 2.160 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.465 2.380 1.030 2.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.720 2.890 3.245 3.400 ;
        RECT  3.015 0.860 3.245 3.400 ;
        RECT  0.900 0.860 3.245 1.200 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.430 3.380 0.770 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.825 -0.180 2.995 0.460 ;
        RECT  0.180 -0.180 0.520 1.200 ;
        END
    END VSS
END NOR4_X0_18_SVT_WB

MACRO NOR3_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR3_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.250 1.620 8.060 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.680 2.330 5.470 2.560 ;
        RECT  5.130 1.915 5.470 2.560 ;
        RECT  0.680 2.220 3.420 2.560 ;
        RECT  2.610 1.915 3.420 2.560 ;
        RECT  0.680 1.760 1.020 2.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.850 1.455 4.660 2.100 ;
        RECT  1.525 1.455 4.660 1.685 ;
        RECT  1.525 1.455 2.225 1.960 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.644  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.330 0.995 8.060 1.225 ;
        RECT  7.720 0.525 8.060 1.225 ;
        RECT  6.040 2.380 7.780 2.720 ;
        RECT  6.040 1.455 6.670 2.720 ;
        RECT  6.330 0.525 6.670 2.720 ;
        RECT  4.890 1.455 6.670 1.685 ;
        RECT  4.890 0.525 5.230 1.685 ;
        RECT  0.900 0.995 5.230 1.225 ;
        RECT  3.570 0.525 3.910 1.225 ;
        RECT  2.240 0.525 2.580 1.225 ;
        RECT  0.900 0.525 1.240 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  4.130 3.515 4.470 4.100 ;
        RECT  1.660 3.515 2.000 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.440 -0.180 8.780 1.225 ;
        RECT  5.610 -0.180 5.950 1.225 ;
        RECT  0.180 -0.180 0.520 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  8.200 2.530 8.540 3.285 ;
        RECT  0.460 2.950 8.540 3.285 ;
    END
END NOR3_X8_18_SVT_WB

MACRO NOR3_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR3_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.505 1.820 6.070 2.205 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.770 1.455 4.340 2.150 ;
        RECT  1.750 1.455 4.340 1.685 ;
        RECT  1.750 1.455 2.090 1.905 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.135 3.330 2.365 ;
        RECT  2.990 1.915 3.330 2.365 ;
        RECT  0.650 1.820 1.030 2.365 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.945  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 2.435 6.540 3.190 ;
        RECT  0.900 0.995 6.540 1.225 ;
        RECT  6.200 0.525 6.540 1.225 ;
        RECT  4.570 2.435 6.540 2.720 ;
        RECT  4.880 0.525 5.220 1.225 ;
        RECT  4.570 0.995 4.920 2.720 ;
        RECT  3.550 0.525 3.890 1.225 ;
        RECT  2.230 0.525 2.570 1.225 ;
        RECT  0.900 0.525 1.240 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  2.770 3.110 3.110 4.100 ;
        RECT  0.180 2.670 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  0.180 -0.180 0.520 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.620 2.595 4.200 2.880 ;
        RECT  3.860 2.595 4.200 3.245 ;
        RECT  3.860 2.950 5.760 3.245 ;
    END
END NOR3_X6_18_SVT_WB

MACRO NOR3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.090 1.670 2.900 2.190 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.420 3.570 2.650 ;
        RECT  3.230 1.860 3.570 2.650 ;
        RECT  1.260 1.770 1.620 2.650 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.210 4.400 1.960 ;
        RECT  0.580 1.210 4.400 1.440 ;
        RECT  0.580 1.210 0.980 1.980 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.320 2.880 4.925 3.220 ;
        RECT  4.630 0.750 4.925 3.220 ;
        RECT  0.785 0.750 4.925 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.310 3.460 4.650 4.100 ;
        RECT  0.320 2.545 0.700 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.080 -0.180 3.420 0.405 ;
        RECT  1.560 -0.180 1.900 0.405 ;
        END
    END VSS
END NOR3_X4_18_SVT_WB

MACRO NOR3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.805 1.535 2.100 2.220 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.620 1.540 2.150 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.580 0.760 2.280 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.623  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.050 2.450 2.620 3.150 ;
        RECT  2.330 0.470 2.620 3.150 ;
        RECT  0.900 0.470 2.620 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.640 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.180 -0.180 0.520 1.350 ;
        END
    END VSS
END NOR3_X2_18_SVT_WB

MACRO NOR3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.595 2.150 2.405 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.175 2.285 1.540 3.115 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.625 1.595 1.030 2.100 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.811  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 0.970 2.660 2.865 ;
        RECT  2.050 2.635 2.390 3.145 ;
        RECT  0.900 0.970 2.660 1.310 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.960 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.660 -0.180 2.470 0.570 ;
        RECT  0.180 -0.180 0.520 1.310 ;
        END
    END VSS
END NOR3_X1_18_SVT_WB

MACRO NOR3_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR3_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.725 1.620 12.230 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.570 1.620 8.080 1.915 ;
        RECT  0.700 2.410 7.800 2.660 ;
        RECT  7.570 1.620 7.800 2.660 ;
        RECT  0.700 2.320 5.860 2.660 ;
        RECT  5.520 1.915 5.860 2.660 ;
        RECT  2.870 2.180 5.860 2.660 ;
        RECT  2.870 1.915 3.210 2.660 ;
        RECT  0.700 1.840 0.930 2.660 ;
        RECT  0.420 1.840 0.930 2.180 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.800 1.455 7.140 2.180 ;
        RECT  1.740 1.455 7.140 1.685 ;
        RECT  4.390 1.455 4.730 1.950 ;
        RECT  1.740 1.455 2.080 1.960 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.966  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 0.885 11.980 1.225 ;
        RECT  11.640 0.525 11.980 1.225 ;
        RECT  8.395 2.475 11.890 2.815 ;
        RECT  10.290 0.525 10.630 1.225 ;
        RECT  8.850 0.525 9.190 1.225 ;
        RECT  8.395 0.885 8.850 2.815 ;
        RECT  7.520 0.525 7.860 1.225 ;
        RECT  6.200 0.525 6.540 1.225 ;
        RECT  4.870 0.525 5.215 1.225 ;
        RECT  3.550 0.525 3.890 1.225 ;
        RECT  2.220 0.525 2.560 1.225 ;
        RECT  0.900 0.525 1.240 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  6.670 3.560 7.010 4.100 ;
        RECT  4.110 3.560 4.450 4.100 ;
        RECT  1.460 3.560 1.800 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  12.360 -0.180 12.700 1.225 ;
        RECT  0.180 -0.180 0.520 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  12.270 2.575 12.610 3.330 ;
        RECT  0.180 3.045 12.610 3.330 ;
        RECT  0.180 3.045 0.520 3.385 ;
    END
END NOR3_X12_18_SVT_WB

MACRO NOR3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.545 2.150 2.355 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 2.330 1.540 2.835 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.395 1.050 2.100 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 0.825 2.660 3.065 ;
        RECT  2.050 2.835 2.390 3.345 ;
        RECT  0.900 0.825 2.660 1.165 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.190 3.350 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.660 -0.180 2.470 0.425 ;
        RECT  0.180 -0.180 0.520 1.165 ;
        END
    END VSS
END NOR3_X0_18_SVT_WB

MACRO NOR2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.850 1.660 4.910 2.100 ;
        RECT  1.230 1.455 4.160 1.685 ;
        RECT  1.230 1.455 2.040 1.915 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.230 2.330 5.565 2.560 ;
        RECT  5.180 1.620 5.565 2.560 ;
        RECT  0.520 2.145 3.470 2.375 ;
        RECT  2.660 1.915 3.470 2.560 ;
        RECT  0.520 1.860 0.860 2.375 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.510  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 2.890 6.025 3.230 ;
        RECT  5.795 0.995 6.025 3.230 ;
        RECT  0.740 0.995 6.025 1.225 ;
        RECT  5.060 0.525 5.400 1.225 ;
        RECT  3.620 0.525 3.960 1.225 ;
        RECT  2.180 0.525 2.520 1.225 ;
        RECT  0.740 0.525 1.080 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.530 3.460 5.870 4.100 ;
        RECT  2.650 3.515 2.990 4.100 ;
        RECT  0.300 2.695 0.640 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.340 -0.180 4.680 0.765 ;
        RECT  2.900 -0.180 3.240 0.765 ;
        RECT  1.460 -0.180 1.800 0.765 ;
        END
    END VSS
END NOR2_X8_18_SVT_WB

MACRO NOR2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.435 1.695 4.300 2.120 ;
        RECT  3.435 1.455 3.675 2.120 ;
        RECT  1.905 1.455 3.675 1.685 ;
        RECT  1.905 1.455 2.245 2.005 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.985 2.235 3.205 2.465 ;
        RECT  2.860 1.915 3.205 2.465 ;
        RECT  0.985 1.770 1.225 2.465 ;
        RECT  0.650 1.770 1.225 2.110 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.138  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.535 0.985 4.825 3.290 ;
        RECT  1.665 2.695 4.825 2.925 ;
        RECT  4.530 0.985 4.825 2.925 ;
        RECT  0.945 0.990 4.825 1.225 ;
        RECT  3.825 0.985 4.825 1.225 ;
        RECT  3.825 0.515 4.165 1.225 ;
        RECT  2.380 0.515 2.725 1.225 ;
        RECT  1.665 2.695 2.005 3.035 ;
        RECT  0.945 0.510 1.285 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.105 3.155 3.445 4.100 ;
        RECT  0.225 2.640 0.565 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.105 -0.180 3.445 0.760 ;
        RECT  1.665 -0.180 2.005 0.760 ;
        END
    END VSS
END NOR2_X6_18_SVT_WB

MACRO NOR2_X5_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.996  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.935 1.595 4.340 1.935 ;
        RECT  1.820 1.595 4.340 1.825 ;
        RECT  1.820 1.595 2.200 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.996  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 3.035 2.870 3.265 ;
        RECT  2.530 2.055 2.870 3.265 ;
        RECT  0.900 2.545 1.130 3.265 ;
        RECT  0.660 2.000 1.030 2.745 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.435  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.110 4.910 2.860 ;
        RECT  0.900 1.110 4.910 1.365 ;
        RECT  0.900 1.055 4.120 1.365 ;
        RECT  3.780 0.540 4.120 1.365 ;
        RECT  2.340 0.540 2.680 1.365 ;
        RECT  1.360 2.520 2.005 2.805 ;
        RECT  1.360 1.055 1.590 2.805 ;
        RECT  0.900 1.055 1.590 1.395 ;
        RECT  0.900 0.540 1.270 1.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.100 2.975 3.400 4.100 ;
        RECT  0.220 2.975 0.505 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.500 -0.180 4.840 0.880 ;
        RECT  3.060 -0.180 3.400 0.825 ;
        RECT  1.620 -0.180 1.960 0.825 ;
        RECT  0.180 -0.180 0.520 1.350 ;
        END
    END VSS
END NOR2_X5_18_SVT_WB

MACRO NOR2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.735 2.120 2.240 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.275 2.785 2.150 ;
        RECT  0.520 1.275 2.785 1.505 ;
        RECT  0.520 1.275 0.860 1.980 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.847  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 2.470 3.245 2.810 ;
        RECT  3.015 0.815 3.245 2.810 ;
        RECT  0.740 0.815 3.245 1.045 ;
        RECT  2.260 0.535 2.660 1.045 ;
        RECT  1.460 2.470 1.800 3.170 ;
        RECT  0.740 0.535 1.080 1.045 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.700 3.105 3.040 4.100 ;
        RECT  0.300 2.635 0.640 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.500 -0.180 1.840 0.405 ;
        END
    END VSS
END NOR2_X4_18_SVT_WB

MACRO NOR2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.320 1.915 2.150 2.660 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.490 1.455 2.785 1.960 ;
        RECT  0.170 1.455 2.785 1.685 ;
        RECT  0.170 1.455 0.980 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.755  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.550 3.070 3.245 3.410 ;
        RECT  3.015 0.470 3.245 3.410 ;
        RECT  2.220 0.470 3.245 1.225 ;
        RECT  0.935 0.470 3.245 0.745 ;
        RECT  0.935 0.470 1.310 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.400 2.380 0.740 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.180 -0.180 0.520 0.875 ;
        END
    END VSS
END NOR2_X3_18_SVT_WB

MACRO NOR2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.175 1.595 1.540 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.480 0.775 2.315 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.159  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.105 2.100 3.300 ;
        RECT  0.960 1.105 2.100 1.335 ;
        RECT  0.960 0.525 1.300 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.175 2.545 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.720 -0.180 2.060 0.875 ;
        RECT  0.240 -0.180 0.580 1.250 ;
        END
    END VSS
END NOR2_X2_18_SVT_WB

MACRO NOR2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.235 1.520 1.575 2.310 ;
        RECT  1.180 1.520 1.575 2.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 2.290 0.980 2.710 ;
        RECT  0.480 1.870 0.820 2.710 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.559  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.680 2.940 2.100 3.280 ;
        RECT  1.805 1.050 2.100 3.280 ;
        RECT  0.960 1.050 2.100 1.280 ;
        RECT  0.960 0.925 1.300 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.195 3.030 0.580 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.720 -0.180 2.060 0.820 ;
        RECT  0.190 -0.180 0.580 1.210 ;
        END
    END VSS
END NOR2_X1_18_SVT_WB

MACRO NOR2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.810 1.710 7.720 2.100 ;
        RECT  6.810 1.455 7.200 2.100 ;
        RECT  1.580 1.455 7.200 1.685 ;
        RECT  3.980 1.455 4.320 2.060 ;
        RECT  1.580 1.455 1.920 2.060 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.980 2.330 8.380 2.715 ;
        RECT  8.040 1.735 8.380 2.715 ;
        RECT  0.760 2.330 8.380 2.560 ;
        RECT  0.760 2.290 5.520 2.560 ;
        RECT  5.180 1.915 5.520 2.560 ;
        RECT  3.020 1.915 3.360 2.560 ;
        RECT  0.760 1.765 1.100 2.560 ;
        RECT  0.260 1.765 1.100 2.105 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.340 2.945 8.845 3.285 ;
        RECT  8.610 0.995 8.845 3.285 ;
        RECT  0.740 0.995 8.845 1.225 ;
        RECT  7.820 0.470 8.160 1.225 ;
        RECT  6.380 0.470 6.720 1.225 ;
        RECT  4.940 0.470 5.280 1.225 ;
        RECT  3.500 0.470 3.840 1.225 ;
        RECT  2.060 0.470 2.400 1.225 ;
        RECT  0.740 0.500 1.080 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.290 3.515 8.630 4.100 ;
        RECT  5.620 3.515 5.960 4.100 ;
        RECT  2.820 3.515 3.160 4.100 ;
        RECT  0.190 2.530 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  7.100 -0.180 7.440 0.760 ;
        RECT  5.660 -0.180 6.000 0.760 ;
        RECT  4.220 -0.180 4.560 0.765 ;
        RECT  2.780 -0.180 3.120 0.765 ;
        END
    END VSS
END NOR2_X12_18_SVT_WB

MACRO NOR2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.195 1.890 1.540 2.805 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.985 0.855 2.860 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.680 3.040 2.100 3.380 ;
        RECT  1.770 1.105 2.100 3.380 ;
        RECT  0.960 1.105 2.100 1.400 ;
        RECT  0.960 1.060 1.300 1.400 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.190 3.095 0.580 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.720 -0.180 2.060 0.875 ;
        RECT  0.190 -0.180 0.580 1.345 ;
        END
    END VSS
END NOR2_X0_18_SVT_WB

MACRO NOR2_A_NOR2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NOR2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.810 2.040 2.150 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 2.380 2.740 2.720 ;
        RECT  2.400 1.840 2.740 2.720 ;
        RECT  0.520 1.675 0.860 2.720 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.680 1.620 7.650 1.960 ;
        RECT  6.680 1.105 6.935 1.960 ;
        RECT  4.450 1.105 6.935 1.390 ;
        RECT  3.980 1.820 4.790 2.180 ;
        RECT  4.450 1.105 4.790 2.180 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.602  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.220 2.940 8.845 3.280 ;
        RECT  8.615 0.580 8.845 3.280 ;
        RECT  3.500 0.580 8.845 0.875 ;
        RECT  3.500 0.470 3.840 0.875 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.350 3.510 8.690 4.100 ;
        RECT  0.310 3.110 0.650 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  7.120 -0.180 7.460 0.350 ;
        RECT  1.460 -0.180 1.800 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 1.105 3.600 1.440 ;
        RECT  5.880 1.620 6.220 2.710 ;
        RECT  5.880 2.370 8.385 2.710 ;
        RECT  8.070 1.840 8.385 2.710 ;
        RECT  3.260 2.410 8.385 2.710 ;
        RECT  3.260 1.105 3.600 3.450 ;
        RECT  1.460 3.110 3.600 3.450 ;
    END
END NOR2_A_NOR2_X8_18_SVT_WB

MACRO NOR2_A_NOR2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NOR2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.680 1.020 2.205 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.250 2.330 1.720 2.765 ;
        RECT  1.380 1.840 1.720 2.765 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.740 1.670 3.275 2.185 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.839  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.220 2.415 4.880 2.755 ;
        RECT  4.650 0.640 4.880 2.755 ;
        RECT  2.420 0.640 4.880 0.980 ;
        RECT  3.220 2.415 3.560 3.225 ;
        RECT  2.420 0.535 2.760 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.390 3.110 4.710 4.100 ;
        RECT  1.660 3.515 2.000 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.660 -0.180 2.000 0.390 ;
        RECT  0.180 -0.180 0.520 1.345 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.535 1.240 1.440 ;
        RECT  0.900 1.210 3.890 1.440 ;
        RECT  3.620 1.210 3.890 1.960 ;
        RECT  3.620 1.620 4.420 1.960 ;
        RECT  2.180 1.210 2.510 3.285 ;
        RECT  0.180 2.995 2.510 3.285 ;
    END
END NOR2_A_NOR2_X4_18_SVT_WB

MACRO NOR2_A_NOR2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NOR2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.750 0.760 2.170 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.095 1.540 1.590 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.790 1.050 3.220 1.695 ;
        RECT  2.790 1.050 3.115 2.080 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.119  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.825 2.380 3.180 3.190 ;
        RECT  2.255 2.380 3.180 2.755 ;
        RECT  2.255 0.630 2.560 2.755 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.460 3.045 1.800 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.180 -0.180 0.520 0.915 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.525 2.025 0.865 ;
        RECT  1.770 0.525 2.025 2.720 ;
        RECT  0.180 2.425 2.025 2.720 ;
    END
END NOR2_A_NOR2_X2_18_SVT_WB

MACRO NOR2_A_NOR2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NOR2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.820 1.030 2.100 ;
        RECT  0.520 1.640 0.860 2.100 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.105 1.560 1.640 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.210 2.785 1.710 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.559  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.690 2.270 3.245 2.735 ;
        RECT  3.015 0.590 3.245 2.735 ;
        RECT  2.315 0.590 3.245 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.500 3.045 1.840 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.220 -0.180 0.475 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.535 2.085 0.875 ;
        RECT  1.790 0.535 2.085 2.720 ;
        RECT  0.310 2.380 2.085 2.720 ;
    END
END NOR2_A_NOR2_X1_18_SVT_WB

MACRO NOR2_A_NOR2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NOR2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.820 1.030 2.100 ;
        RECT  0.420 1.540 0.760 2.100 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.070 1.540 1.605 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 1.700 2.680 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.480 2.420 3.245 2.760 ;
        RECT  2.910 0.500 3.245 2.760 ;
        RECT  2.230 0.500 3.245 0.840 ;
        RECT  2.480 2.420 2.820 3.205 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.330 2.865 1.670 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.180 -0.180 0.520 0.840 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.500 2.000 0.840 ;
        RECT  1.770 1.070 2.150 1.410 ;
        RECT  1.770 0.500 2.000 2.635 ;
        RECT  0.180 2.330 2.000 2.635 ;
        RECT  0.180 2.330 0.520 3.205 ;
    END
END NOR2_A_NOR2_X0_18_SVT_WB

MACRO NOR2_A_NAND3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NAND3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.770 1.540 2.275 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.260 1.030 1.560 ;
        RECT  0.420 1.260 0.760 1.960 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.785 2.135 4.900 2.365 ;
        RECT  4.560 1.915 4.900 2.365 ;
        RECT  2.785 1.770 3.220 2.365 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.455 4.900 1.685 ;
        RECT  4.560 1.210 4.900 1.685 ;
        RECT  3.450 1.455 3.790 1.905 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.603  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 2.595 5.510 2.935 ;
        RECT  5.130 2.380 5.510 2.935 ;
        RECT  2.800 0.940 3.980 1.225 ;
        RECT  2.325 1.225 3.140 1.525 ;
        RECT  2.325 1.225 2.555 2.935 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.360 3.165 4.700 4.100 ;
        RECT  2.920 3.165 3.260 4.100 ;
        RECT  1.330 3.110 1.670 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  5.685 -0.180 5.970 1.410 ;
        RECT  1.660 -0.180 2.000 0.405 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.535 1.240 0.875 ;
        RECT  2.230 0.410 5.360 0.710 ;
        RECT  0.900 0.635 2.570 0.875 ;
        RECT  5.130 0.410 5.360 1.980 ;
        RECT  1.770 0.635 2.095 1.960 ;
        RECT  5.130 1.640 5.635 1.980 ;
        RECT  1.770 0.635 2.000 2.880 ;
        RECT  0.180 2.540 2.000 2.880 ;
        RECT  0.180 2.380 0.520 3.190 ;
    END
END NOR2_A_NAND3_X4_18_SVT_WB

MACRO NOR2_A_NAND3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NAND3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.200 1.385 1.540 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.770 0.915 2.150 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.930 0.850 3.270 1.965 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.625 3.885 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.677  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.840 2.420 4.345 3.230 ;
        RECT  4.115 0.480 4.345 3.230 ;
        RECT  3.840 0.480 4.345 1.395 ;
        RECT  2.450 2.420 4.345 2.760 ;
        RECT  2.450 2.420 2.790 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.170 3.110 3.510 4.100 ;
        RECT  1.730 3.110 2.070 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  2.075 -0.180 2.360 0.810 ;
        RECT  0.190 -0.180 0.530 0.915 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.910 0.575 1.845 0.915 ;
        RECT  1.615 0.575 1.845 2.720 ;
        RECT  1.615 1.845 2.570 2.185 ;
        RECT  1.615 1.845 1.955 2.720 ;
        RECT  0.190 2.380 1.955 2.720 ;
    END
END NOR2_A_NAND3_X2_18_SVT_WB

MACRO NOR2_A_NAND3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NAND3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.070 1.590 1.540 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.820 1.030 2.100 ;
        RECT  0.420 1.540 0.760 2.100 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 1.820 2.710 2.355 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.515 3.260 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.839  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.050 2.790 3.780 3.115 ;
        RECT  3.490 0.615 3.780 3.115 ;
        RECT  3.200 0.825 3.780 1.165 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.365 3.515 2.980 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.180 -0.180 0.520 0.840 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.500 2.160 0.840 ;
        RECT  1.820 0.500 2.160 1.630 ;
        RECT  1.820 0.500 2.070 2.560 ;
        RECT  0.180 2.330 2.070 2.560 ;
        RECT  0.180 2.330 0.520 2.960 ;
    END
END NOR2_A_NAND3_X1_18_SVT_WB

MACRO NOR2_A_NAND3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_NAND3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.070 1.400 1.395 1.800 ;
        RECT  0.135 1.400 1.395 1.645 ;
        RECT  0.135 1.115 0.550 1.645 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.250 2.335 1.060 2.670 ;
        RECT  0.250 2.055 0.745 2.670 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 2.255 2.935 2.530 ;
        RECT  2.330 1.640 2.660 2.530 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.260 3.270 1.955 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.065 2.775 3.780 3.115 ;
        RECT  3.505 0.665 3.780 3.115 ;
        RECT  3.370 2.170 3.780 3.115 ;
        RECT  3.455 0.665 3.780 1.075 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.370 3.515 2.985 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.175 -0.180 1.915 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.860 0.860 1.885 1.145 ;
        RECT  1.625 0.860 1.885 2.530 ;
        RECT  1.510 2.205 1.835 3.275 ;
        RECT  0.180 2.995 1.835 3.275 ;
    END
END NOR2_A_NAND3_X0_18_SVT_WB

MACRO NOR2_A_AOI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_AOI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.760 0.735 2.150 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.975 1.095 1.540 1.905 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.520 1.260 2.805 1.980 ;
        RECT  2.300 1.260 2.805 1.600 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.495 1.765 3.825 2.380 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.150 2.695 8.010 3.265 ;
        RECT  7.180 2.565 8.010 3.265 ;
        RECT  7.180 1.080 8.010 1.420 ;
        RECT  7.670 0.675 8.010 1.420 ;
        RECT  7.180 1.080 7.560 3.265 ;
        RECT  6.150 1.080 8.010 1.345 ;
        RECT  6.150 2.695 6.490 3.450 ;
        RECT  6.150 0.540 6.490 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.390 2.565 8.730 4.100 ;
        RECT  6.910 3.510 7.250 4.100 ;
        RECT  5.390 3.515 5.730 4.100 ;
        RECT  0.780 3.515 1.590 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.390 -0.180 8.730 1.375 ;
        RECT  6.910 -0.180 7.250 0.850 ;
        RECT  5.390 -0.180 5.730 0.405 ;
        RECT  3.790 -0.180 4.130 0.400 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.860 0.470 2.070 0.810 ;
        RECT  1.770 0.470 2.070 2.335 ;
        RECT  1.540 2.140 1.905 2.740 ;
        RECT  0.190 2.380 1.905 2.740 ;
        RECT  2.010 3.045 3.790 3.385 ;
        RECT  2.300 0.630 4.640 0.915 ;
        RECT  4.410 0.630 4.640 1.980 ;
        RECT  4.410 1.640 4.875 1.980 ;
        RECT  3.035 0.630 3.265 2.720 ;
        RECT  2.730 2.370 3.265 2.720 ;
        RECT  4.870 0.805 5.335 1.145 ;
        RECT  5.105 1.620 6.665 1.960 ;
        RECT  5.105 0.805 5.335 2.720 ;
        RECT  4.830 2.380 5.335 2.720 ;
    END
END NOR2_A_AOI21_X8_18_SVT_WB

MACRO NOR2_A_AOI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_AOI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.485 1.820 1.030 2.100 ;
        RECT  0.485 1.590 0.825 2.100 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.450 1.595 2.150 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.495 1.820 4.950 2.200 ;
        RECT  2.850 2.135 4.720 2.365 ;
        RECT  2.850 1.860 3.135 2.365 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.260 3.830 1.905 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.628  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.390 2.595 5.545 2.880 ;
        RECT  5.180 2.330 5.545 2.880 ;
        RECT  5.180 1.100 5.430 2.880 ;
        RECT  2.390 1.100 2.825 1.440 ;
        RECT  2.390 1.100 2.620 2.880 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  5.865 2.640 6.205 4.100 ;
        RECT  1.545 3.110 1.885 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.140 -0.180 6.445 1.280 ;
        RECT  3.715 -0.180 4.055 0.405 ;
        RECT  1.725 -0.180 2.065 0.405 ;
        RECT  0.245 -0.180 0.585 1.345 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.265 3.110 5.485 3.450 ;
        RECT  0.965 0.535 1.305 0.875 ;
        RECT  0.965 0.635 5.910 0.870 ;
        RECT  0.965 0.635 2.160 0.875 ;
        RECT  5.660 0.635 5.910 1.960 ;
        RECT  1.875 0.635 2.160 2.720 ;
        RECT  0.245 2.380 2.160 2.720 ;
        RECT  0.245 2.380 0.585 3.190 ;
    END
END NOR2_A_AOI21_X4_18_SVT_WB

MACRO NOR2_A_AOI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_AOI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.090 0.760 2.425 ;
        RECT  0.140 1.715 0.490 2.425 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.980 1.210 1.545 1.660 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.430 1.260 2.710 1.960 ;
        RECT  2.255 1.260 2.710 1.600 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.555 3.780 2.245 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.650 2.380 3.220 2.720 ;
        RECT  2.940 0.640 3.220 2.720 ;
        RECT  2.245 0.640 3.220 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.165 3.515 1.515 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.390 -0.180 3.730 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.690 2.015 0.980 ;
        RECT  1.275 2.490 2.015 2.730 ;
        RECT  1.775 0.690 2.015 2.730 ;
        RECT  0.180 2.705 1.505 3.065 ;
        RECT  1.930 3.045 3.710 3.385 ;
    END
END NOR2_A_AOI21_X2_18_SVT_WB

MACRO NOR2_A_AOI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_AOI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.415 1.190 0.980 1.590 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.955 1.540 2.235 ;
        RECT  1.210 1.660 1.540 2.235 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.255 1.880 2.705 2.200 ;
        RECT  2.365 1.660 2.705 2.200 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.495 3.780 2.150 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.760 2.430 3.220 2.770 ;
        RECT  2.935 0.620 3.220 2.770 ;
        RECT  2.385 0.620 3.220 0.960 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.400 3.515 1.740 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.170 -0.180 0.535 0.960 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.620 2.155 0.960 ;
        RECT  1.795 0.620 2.155 1.530 ;
        RECT  1.795 0.620 2.025 3.005 ;
        RECT  0.175 2.720 2.025 3.005 ;
        RECT  0.175 2.720 0.610 3.060 ;
    END
END NOR2_A_AOI21_X1_18_SVT_WB

MACRO NOR2_A_AOI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2_A_AOI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.425 1.190 0.980 1.590 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.010 1.955 1.540 2.235 ;
        RECT  1.210 1.660 1.540 2.235 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.870 2.710 2.150 ;
        RECT  2.365 1.555 2.710 2.150 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 0.935 3.780 1.590 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.760 2.380 3.220 2.720 ;
        RECT  2.940 0.590 3.220 2.720 ;
        RECT  2.370 0.590 3.220 0.930 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.330 3.515 1.670 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.220 -0.180 0.480 0.940 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.590 1.280 0.960 ;
        RECT  0.940 0.730 2.140 0.960 ;
        RECT  1.800 0.730 2.140 1.450 ;
        RECT  1.800 0.730 2.030 2.970 ;
        RECT  0.180 2.630 2.030 2.970 ;
    END
END NOR2_A_AOI21_X0_18_SVT_WB

MACRO NOR2P3_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.015 1.065 6.580 1.885 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.635 0.740 1.930 ;
        RECT  0.140 1.165 0.685 1.930 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.888  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.050 5.785 1.280 ;
        RECT  5.460 0.535 5.785 1.280 ;
        RECT  5.380 1.765 5.720 3.035 ;
        RECT  3.940 1.765 5.720 1.995 ;
        RECT  3.940 0.535 4.280 2.815 ;
        RECT  2.380 0.535 2.760 1.280 ;
        RECT  0.915 0.535 1.240 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  2.460 2.630 2.800 4.100 ;
        RECT  0.940 2.630 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.180 -0.180 6.520 0.835 ;
        RECT  4.700 -0.180 5.040 0.820 ;
        RECT  3.180 -0.180 3.520 0.820 ;
        RECT  1.660 -0.180 2.000 0.820 ;
        RECT  0.180 -0.180 0.520 0.835 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.160 3.560 2.400 ;
        RECT  0.180 2.160 0.520 3.135 ;
        RECT  3.220 2.160 3.560 3.505 ;
        RECT  4.660 2.225 5.000 3.505 ;
        RECT  3.220 3.165 5.000 3.505 ;
        RECT  1.700 2.160 2.040 3.330 ;
        RECT  6.140 2.695 6.480 3.505 ;
        RECT  3.220 3.265 6.480 3.505 ;
    END
END NOR2P3_X8_18_SVT_WB

MACRO NOR2P3_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.075  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.065 4.435 1.605 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.075  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.070 0.680 1.880 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.258  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.500 2.115 4.840 3.285 ;
        RECT  3.060 2.115 4.840 2.400 ;
        RECT  3.600 0.470 4.120 0.810 ;
        RECT  3.060 1.025 3.830 2.400 ;
        RECT  3.600 0.470 3.830 2.400 ;
        RECT  0.910 1.025 3.830 1.255 ;
        RECT  2.340 0.470 2.680 1.255 ;
        RECT  0.910 0.470 1.240 1.255 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  1.620 2.685 1.960 4.100 ;
        RECT  0.180 2.640 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.500 -0.180 4.840 0.810 ;
        RECT  3.060 -0.180 3.370 0.795 ;
        RECT  1.620 -0.180 1.960 0.795 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.225 2.680 2.455 ;
        RECT  2.340 2.225 2.680 3.450 ;
        RECT  0.900 2.225 1.240 3.450 ;
        RECT  2.340 2.640 4.120 3.450 ;
    END
END NOR2P3_X6_18_SVT_WB

MACRO NOR2P3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.648  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.985 1.210 3.780 1.975 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.648  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.240 1.460 1.580 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.345  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.465 0.670 2.755 2.790 ;
        RECT  0.945 0.670 2.755 1.010 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.985 2.630 1.325 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.205 -0.180 3.545 0.955 ;
        RECT  1.705 -0.180 2.045 0.440 ;
        RECT  0.175 -0.180 0.565 0.955 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.225 2.170 2.085 2.400 ;
        RECT  1.745 2.170 2.085 3.385 ;
        RECT  0.225 2.170 0.565 3.330 ;
        RECT  3.225 2.505 3.565 3.385 ;
        RECT  1.745 3.045 3.565 3.385 ;
    END
END NOR2P3_X4_18_SVT_WB

MACRO NOR2P3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.215 1.390 1.540 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.445 0.525 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.779  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.435 1.720 3.220 ;
        RECT  0.755 0.870 1.280 1.160 ;
        RECT  0.755 2.435 1.720 2.775 ;
        RECT  0.755 0.870 0.985 2.775 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.175 2.380 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.700 -0.180 2.040 0.890 ;
        RECT  0.180 -0.180 0.520 0.890 ;
        END
    END VSS
END NOR2P3_X2_18_SVT_WB

MACRO NOR2P3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.205 1.530 1.545 2.285 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.158  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.585 0.515 2.285 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.537  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.745 2.520 1.710 3.220 ;
        RECT  0.745 1.050 1.320 1.300 ;
        RECT  0.745 1.050 0.975 3.220 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.180 2.520 0.515 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.180 -0.180 1.955 0.820 ;
        END
    END VSS
END NOR2P3_X1_18_SVT_WB

MACRO NOR2P3_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.065  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.900 1.170 12.240 1.930 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.065  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.430 0.835 2.195 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.166  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.655 0.600 12.515 0.940 ;
        RECT  11.375 2.075 11.715 2.915 ;
        RECT  0.255 0.970 11.455 1.200 ;
        RECT  10.655 0.600 11.455 1.200 ;
        RECT  7.055 2.075 11.715 2.345 ;
        RECT  9.935 2.075 10.275 2.915 ;
        RECT  9.085 0.970 9.565 2.345 ;
        RECT  3.135 0.860 9.555 1.200 ;
        RECT  9.215 0.535 9.555 2.345 ;
        RECT  8.495 2.075 8.835 2.915 ;
        RECT  7.695 0.535 8.035 1.200 ;
        RECT  7.055 2.075 7.395 2.915 ;
        RECT  4.655 0.850 6.515 1.200 ;
        RECT  6.175 0.535 6.515 1.200 ;
        RECT  4.655 0.535 4.995 1.200 ;
        RECT  3.135 0.535 3.475 1.200 ;
        RECT  1.695 0.600 2.035 1.200 ;
        RECT  0.255 0.600 0.595 1.200 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  5.575 3.045 5.915 4.100 ;
        RECT  4.055 3.045 4.395 4.100 ;
        RECT  2.535 3.045 2.875 4.100 ;
        RECT  1.015 3.045 1.355 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  11.415 -0.180 11.755 0.370 ;
        RECT  9.935 -0.180 10.275 0.740 ;
        RECT  8.455 -0.180 8.795 0.405 ;
        RECT  6.935 -0.180 7.275 0.405 ;
        RECT  5.415 -0.180 5.755 0.405 ;
        RECT  3.895 -0.180 4.235 0.405 ;
        RECT  2.415 -0.180 2.755 0.740 ;
        RECT  0.975 -0.180 1.315 0.740 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.255 2.575 6.675 2.815 ;
        RECT  6.335 2.575 6.675 3.385 ;
        RECT  7.775 2.575 8.115 3.385 ;
        RECT  9.215 2.575 9.555 3.385 ;
        RECT  10.655 2.575 10.995 3.385 ;
        RECT  0.255 2.575 0.595 3.385 ;
        RECT  1.775 2.575 2.115 3.385 ;
        RECT  3.295 2.575 3.635 3.385 ;
        RECT  4.815 2.575 5.155 3.385 ;
        RECT  12.135 2.530 12.475 3.385 ;
        RECT  6.335 3.145 12.475 3.385 ;
    END
END NOR2P3_X16_18_SVT_WB

MACRO NOR2P3_X14_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3_X14_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.682  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.440 1.200 11.060 1.995 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.682  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.445 0.790 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.304  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.680 2.225 11.020 3.145 ;
        RECT  7.800 2.225 11.020 2.465 ;
        RECT  0.940 0.970 10.210 1.200 ;
        RECT  9.900 0.600 10.210 1.200 ;
        RECT  9.240 2.225 9.580 2.925 ;
        RECT  2.380 0.860 8.800 1.200 ;
        RECT  8.460 0.535 8.800 1.200 ;
        RECT  7.800 0.860 8.185 2.465 ;
        RECT  7.800 0.860 8.140 2.925 ;
        RECT  6.360 0.860 8.185 2.100 ;
        RECT  6.940 0.535 7.280 2.100 ;
        RECT  6.360 0.860 6.700 2.925 ;
        RECT  5.420 0.535 5.760 1.200 ;
        RECT  3.900 0.535 4.240 1.200 ;
        RECT  2.380 0.535 2.720 1.200 ;
        RECT  0.940 0.600 1.280 1.200 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  4.880 3.100 5.220 4.100 ;
        RECT  3.360 3.100 3.700 4.100 ;
        RECT  1.840 3.100 2.180 4.100 ;
        RECT  0.360 2.515 0.700 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  10.660 -0.180 11.000 0.470 ;
        RECT  9.180 -0.180 9.520 0.740 ;
        RECT  7.700 -0.180 8.040 0.405 ;
        RECT  6.180 -0.180 6.520 0.405 ;
        RECT  4.660 -0.180 5.000 0.405 ;
        RECT  3.140 -0.180 3.480 0.405 ;
        RECT  1.660 -0.180 2.000 0.740 ;
        RECT  0.180 -0.180 0.520 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.080 2.410 5.980 2.750 ;
        RECT  2.600 2.410 4.460 2.825 ;
        RECT  2.600 2.410 2.940 3.110 ;
        RECT  5.640 2.410 5.980 3.450 ;
        RECT  7.080 2.695 7.420 3.450 ;
        RECT  8.520 2.695 8.860 3.450 ;
        RECT  1.080 2.410 1.420 3.275 ;
        RECT  4.120 2.410 4.460 3.330 ;
        RECT  9.960 2.695 10.300 3.450 ;
        RECT  5.640 3.155 10.300 3.450 ;
    END
END NOR2P3_X14_18_SVT_WB

MACRO NOR2P3T_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3T_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.075  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.415 1.375 6.030 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.463  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.580 0.975 1.875 ;
        RECT  0.140 1.165 0.515 1.875 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.498  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.595 2.525 5.935 3.280 ;
        RECT  5.595 0.550 5.915 1.115 ;
        RECT  4.010 2.525 5.935 2.765 ;
        RECT  4.055 0.885 5.915 1.115 ;
        RECT  4.010 1.050 4.495 2.765 ;
        RECT  4.055 0.535 4.435 2.765 ;
        RECT  1.015 1.050 4.495 1.280 ;
        RECT  2.535 0.535 2.875 1.280 ;
        RECT  1.015 0.535 1.355 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  2.675 2.630 3.015 4.100 ;
        RECT  1.155 2.575 1.495 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.815 -0.180 5.155 0.655 ;
        RECT  3.295 -0.180 3.635 0.820 ;
        RECT  1.775 -0.180 2.115 0.820 ;
        RECT  0.255 -0.180 0.595 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.395 2.105 3.775 2.345 ;
        RECT  1.915 2.105 3.775 2.400 ;
        RECT  3.435 2.105 3.775 3.500 ;
        RECT  0.395 2.105 0.735 3.275 ;
        RECT  1.915 2.105 2.255 3.275 ;
        RECT  3.435 2.995 5.215 3.500 ;
    END
END NOR2P3T_X6_18_SVT_WB

MACRO NOR2P3T_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3T_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.671  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.750 1.445 4.355 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.046  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.125 0.760 1.935 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.653  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.900 0.550 4.240 1.215 ;
        RECT  2.380 0.985 4.240 1.215 ;
        RECT  3.180 0.985 3.520 3.035 ;
        RECT  0.990 1.065 3.520 1.295 ;
        RECT  2.380 0.550 2.800 1.295 ;
        RECT  0.990 0.550 1.280 1.295 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  1.700 2.555 2.040 4.100 ;
        RECT  0.220 2.555 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.180 -0.180 3.520 0.755 ;
        RECT  1.700 -0.180 2.040 0.835 ;
        RECT  0.220 -0.180 0.560 0.835 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 2.085 2.800 2.325 ;
        RECT  0.940 2.085 1.280 3.255 ;
        RECT  2.460 2.085 2.800 3.505 ;
        RECT  3.940 2.555 4.280 3.505 ;
        RECT  2.460 3.265 4.280 3.505 ;
    END
END NOR2P3T_X4_18_SVT_WB

MACRO NOR2P3T_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3T_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.335 1.390 2.660 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.648  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.210 1.480 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.011  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.525 2.585 3.120 2.925 ;
        RECT  2.890 0.670 3.120 2.925 ;
        RECT  0.965 0.670 3.120 0.980 ;
        RECT  2.525 2.585 2.865 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.005 3.100 1.345 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.725 -0.180 2.065 0.440 ;
        RECT  0.245 -0.180 0.585 0.955 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.245 2.115 2.105 2.455 ;
        RECT  1.765 2.115 2.105 3.285 ;
        RECT  0.245 2.115 0.585 3.330 ;
    END
END NOR2P3T_X2_18_SVT_WB

MACRO NOR2P3T_X10_18_SVT_WB
    CLASS CORE ;
    FOREIGN NOR2P3T_X10_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.890  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.320 1.120 9.940 1.885 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.682  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.175 0.780 1.930 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.139  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.540 2.115 9.880 3.135 ;
        RECT  6.640 2.115 9.880 2.425 ;
        RECT  1.195 1.105 9.090 1.335 ;
        RECT  8.800 0.470 9.090 1.335 ;
        RECT  8.080 2.115 8.420 2.885 ;
        RECT  7.280 0.470 7.620 1.335 ;
        RECT  6.640 1.105 7.140 2.425 ;
        RECT  6.640 1.105 6.980 2.870 ;
        RECT  2.715 1.050 6.100 1.335 ;
        RECT  5.760 0.470 6.100 1.335 ;
        RECT  2.715 0.970 4.575 1.335 ;
        RECT  4.235 0.535 4.575 1.335 ;
        RECT  2.715 0.535 3.055 1.335 ;
        RECT  1.195 0.600 1.535 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  4.775 2.630 5.115 4.100 ;
        RECT  3.295 2.630 3.635 4.100 ;
        RECT  1.815 2.710 2.155 4.100 ;
        RECT  0.375 2.575 0.715 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  9.560 -0.180 9.900 0.890 ;
        RECT  8.040 -0.180 8.380 0.875 ;
        RECT  6.520 -0.180 6.860 0.875 ;
        RECT  4.995 -0.180 5.335 0.820 ;
        RECT  3.475 -0.180 3.815 0.405 ;
        RECT  1.955 -0.180 2.295 0.875 ;
        RECT  0.435 -0.180 0.775 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.095 2.060 5.915 2.400 ;
        RECT  1.095 2.060 2.875 2.410 ;
        RECT  5.575 2.060 5.915 3.410 ;
        RECT  7.360 2.655 7.700 3.410 ;
        RECT  5.575 3.100 7.700 3.410 ;
        RECT  1.095 2.060 1.435 3.190 ;
        RECT  2.535 2.060 2.875 3.330 ;
        RECT  4.055 2.060 4.395 3.330 ;
        RECT  8.800 2.655 9.140 3.410 ;
        RECT  5.575 3.115 9.140 3.410 ;
    END
END NOR2P3T_X10_18_SVT_WB

MACRO NAND4_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.540 2.330 10.020 2.660 ;
        RECT  9.680 1.915 10.020 2.660 ;
        RECT  7.540 1.915 7.880 2.660 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.740 1.455 11.080 1.960 ;
        RECT  6.210 1.455 11.080 1.685 ;
        RECT  8.240 1.455 9.050 2.100 ;
        RECT  6.210 1.455 6.550 1.980 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.180 1.360 5.550 2.200 ;
        RECT  2.710 1.360 5.550 1.630 ;
        RECT  2.710 1.360 3.520 1.905 ;
        RECT  0.765 1.360 5.550 1.590 ;
        RECT  0.765 1.360 1.050 1.960 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.380 2.135 4.230 2.365 ;
        RECT  3.890 1.860 4.230 2.365 ;
        RECT  1.380 1.820 2.190 2.365 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.165  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.800 2.190 11.645 2.425 ;
        RECT  11.310 0.985 11.645 2.425 ;
        RECT  7.330 0.985 11.645 1.225 ;
        RECT  6.430 3.110 11.030 3.450 ;
        RECT  10.800 2.190 11.030 3.450 ;
        RECT  10.520 2.640 11.030 3.450 ;
        RECT  6.430 2.640 6.770 3.450 ;
        RECT  0.900 2.640 6.770 2.950 ;
        RECT  4.990 2.640 5.330 3.450 ;
        RECT  3.670 2.640 4.010 3.450 ;
        RECT  2.230 2.640 2.570 3.450 ;
        RECT  0.900 2.640 1.240 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  11.260 2.655 11.580 4.100 ;
        RECT  5.710 3.180 6.050 4.100 ;
        RECT  0.180 2.655 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  4.140 -0.180 4.480 0.405 ;
        RECT  1.660 -0.180 2.000 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.250 0.535 0.590 0.975 ;
        RECT  4.705 0.470 11.300 0.755 ;
        RECT  0.250 0.635 5.045 0.975 ;
        RECT  0.250 0.535 0.535 1.345 ;
    END
END NAND4_X8_18_SVT_WB

MACRO NAND4_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.940 1.455 8.260 2.150 ;
        RECT  5.910 1.455 8.260 1.685 ;
        RECT  5.910 1.455 6.250 1.905 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.570 2.135 7.380 2.365 ;
        RECT  7.040 1.915 7.380 2.365 ;
        RECT  4.570 1.820 4.950 2.365 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.135 4.340 2.365 ;
        RECT  3.870 1.770 4.340 2.365 ;
        RECT  1.740 1.910 2.080 2.365 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.970 1.450 3.310 1.905 ;
        RECT  0.420 1.450 3.310 1.680 ;
        RECT  0.420 1.450 0.980 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.860  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.655 8.820 2.950 ;
        RECT  8.490 0.605 8.820 2.950 ;
        RECT  5.670 0.995 8.820 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.440 3.180 8.780 4.100 ;
        RECT  4.350 3.180 4.690 4.100 ;
        RECT  0.180 2.635 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  2.690 -0.180 3.030 0.405 ;
        RECT  0.180 -0.180 0.520 0.795 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.255 0.470 7.160 0.765 ;
        RECT  3.255 0.470 3.595 1.220 ;
        RECT  1.500 0.925 3.595 1.220 ;
    END
END NAND4_X6_18_SVT_WB

MACRO NAND4_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.490 1.450 5.460 1.680 ;
        RECT  5.120 1.210 5.460 1.680 ;
        RECT  4.490 1.450 4.830 1.960 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.480 2.190 5.550 2.420 ;
        RECT  5.210 1.910 5.550 2.420 ;
        RECT  3.480 1.770 3.780 2.420 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 2.135 2.790 2.365 ;
        RECT  2.505 1.860 2.790 2.365 ;
        RECT  0.660 1.770 1.000 2.365 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.210 1.720 1.905 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.051  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.695 5.310 3.395 ;
        RECT  3.020 0.935 4.660 1.220 ;
        RECT  3.020 0.935 3.250 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  0.180 2.695 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  1.590 -0.180 1.930 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.150 0.475 5.975 0.705 ;
        RECT  0.400 0.635 2.490 0.975 ;
        RECT  0.400 0.635 0.740 1.335 ;
        RECT  5.690 0.475 5.975 1.440 ;
    END
END NAND4_X4_18_SVT_WB

MACRO NAND4_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.265 2.320 2.780 2.660 ;
        RECT  2.495 1.840 2.780 2.660 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.260 2.395 1.600 ;
        RECT  1.770 1.260 2.165 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.450 1.540 2.150 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.635 0.980 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.746  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.915 3.110 3.240 3.450 ;
        RECT  3.010 0.630 3.240 3.450 ;
        RECT  2.735 0.630 3.240 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.195 2.640 0.535 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.195 -0.180 0.535 1.405 ;
        END
    END VSS
END NAND4_X2_18_SVT_WB

MACRO NAND4_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.505 2.720 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.055 2.100 1.590 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.820 1.590 2.275 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.230 1.230 1.590 ;
        RECT  0.900 1.000 1.230 1.590 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.952  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.775 3.180 3.220 ;
        RECT  2.950 0.710 3.180 3.220 ;
        RECT  2.765 0.710 3.180 1.050 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.660 3.515 3.165 4.100 ;
        RECT  0.180 2.775 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.180 -0.180 0.465 1.000 ;
        END
    END VSS
END NAND4_X1_18_SVT_WB

MACRO NAND4_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.740 1.455 16.150 2.100 ;
        RECT  10.270 1.455 16.150 1.685 ;
        RECT  13.320 1.455 13.660 1.915 ;
        RECT  10.270 1.455 10.610 1.915 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.500 1.620 17.240 1.915 ;
        RECT  14.560 2.330 16.730 2.660 ;
        RECT  16.500 1.620 16.730 2.660 ;
        RECT  9.240 2.145 14.790 2.375 ;
        RECT  14.280 1.915 14.790 2.375 ;
        RECT  11.400 1.915 11.740 2.375 ;
        RECT  9.240 1.860 9.580 2.375 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.280 1.455 8.620 1.980 ;
        RECT  0.650 1.455 8.620 1.685 ;
        RECT  6.120 1.455 6.460 1.915 ;
        RECT  2.840 1.455 3.180 1.915 ;
        RECT  0.650 1.455 1.030 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.145 7.420 2.375 ;
        RECT  7.080 1.915 7.420 2.375 ;
        RECT  4.260 1.915 4.600 2.375 ;
        RECT  1.770 1.915 2.150 2.660 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.342  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.960 2.145 17.805 2.425 ;
        RECT  17.470 0.995 17.805 2.425 ;
        RECT  10.490 0.995 17.805 1.225 ;
        RECT  13.800 3.110 17.190 3.450 ;
        RECT  16.960 2.145 17.190 3.450 ;
        RECT  16.680 2.890 17.190 3.450 ;
        RECT  13.800 2.640 14.140 3.450 ;
        RECT  2.380 2.640 14.140 2.895 ;
        RECT  12.360 2.640 12.700 3.395 ;
        RECT  10.920 2.640 11.260 3.395 ;
        RECT  9.480 2.640 9.820 3.395 ;
        RECT  8.040 2.640 8.380 3.395 ;
        RECT  6.600 2.640 6.940 3.395 ;
        RECT  5.220 2.640 5.560 3.395 ;
        RECT  3.780 2.640 4.120 3.395 ;
        RECT  0.900 2.890 2.680 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  17.420 2.655 17.740 4.100 ;
        RECT  13.080 3.135 13.420 4.100 ;
        RECT  8.760 3.125 9.100 4.100 ;
        RECT  4.500 3.180 4.840 4.100 ;
        RECT  0.180 2.695 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  7.070 -0.180 7.410 0.405 ;
        RECT  4.500 -0.180 4.840 0.740 ;
        RECT  1.760 -0.180 2.100 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  7.815 0.470 17.460 0.765 ;
        RECT  7.815 0.470 8.155 1.225 ;
        RECT  0.460 0.970 8.155 1.225 ;
    END
END NAND4_X12_18_SVT_WB

MACRO NAND4_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.640 2.785 2.175 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 0.650 2.150 1.510 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.125 1.820 1.695 2.210 ;
        RECT  1.125 1.820 1.465 2.490 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.210 1.270 1.590 ;
        RECT  1.040 0.905 1.270 1.590 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.720 3.245 3.060 ;
        RECT  3.015 0.650 3.245 3.060 ;
        RECT  2.720 0.650 3.245 1.030 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.665 3.460 3.170 4.100 ;
        RECT  0.180 2.720 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.470 -0.180 0.810 0.980 ;
        END
    END VSS
END NAND4_X0_18_SVT_WB

MACRO NAND4T_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.110 1.595 16.975 2.145 ;
        RECT  15.110 1.595 15.700 2.275 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.306  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.165 1.750 14.470 2.385 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.369  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.860 1.755 9.145 2.385 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.337  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.065 1.750 4.720 2.385 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.180 2.630 17.720 2.860 ;
        RECT  17.380 1.045 17.720 2.860 ;
        RECT  15.940 2.380 17.720 2.860 ;
        RECT  15.940 1.045 17.720 1.345 ;
        RECT  14.500 2.630 14.840 3.145 ;
        RECT  13.060 2.630 13.400 3.145 ;
        RECT  11.620 2.630 11.960 3.145 ;
        RECT  9.500 2.380 11.765 2.860 ;
        RECT  10.180 2.380 10.520 3.145 ;
        RECT  8.740 2.630 9.080 3.145 ;
        RECT  7.300 2.630 7.640 3.145 ;
        RECT  5.860 2.630 6.200 3.145 ;
        RECT  4.420 2.630 4.760 3.145 ;
        RECT  2.980 2.630 3.320 3.145 ;
        RECT  0.180 2.630 1.880 3.145 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 19.040 4.100 ;
        RECT  18.100 3.110 18.440 4.100 ;
        RECT  16.660 3.160 17.000 4.100 ;
        RECT  15.220 3.090 15.560 4.100 ;
        RECT  13.780 3.095 14.120 4.100 ;
        RECT  12.340 3.095 12.680 4.100 ;
        RECT  10.900 3.090 11.240 4.100 ;
        RECT  9.460 3.090 9.800 4.100 ;
        RECT  8.020 3.090 8.360 4.100 ;
        RECT  6.580 3.090 6.920 4.100 ;
        RECT  5.140 3.090 5.480 4.100 ;
        RECT  3.700 3.090 4.040 4.100 ;
        RECT  2.260 3.090 2.600 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 19.040 0.180 ;
        RECT  4.420 -0.180 4.760 0.770 ;
        RECT  2.980 -0.180 3.320 0.770 ;
        RECT  0.180 -0.180 0.520 0.770 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  5.140 0.470 9.800 0.810 ;
        RECT  5.140 0.470 5.480 1.340 ;
        RECT  0.900 1.000 5.480 1.340 ;
        RECT  5.860 1.040 14.840 1.380 ;
        RECT  10.900 0.470 18.440 0.810 ;
    END
END NAND4T_X8_18_SVT_WB

MACRO NAND4T_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.180 1.620 11.700 2.410 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.709  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.775 1.730 10.645 2.370 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.804  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.715 1.745 7.435 2.375 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.757  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.855 1.760 3.550 2.390 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.345 0.685 13.765 3.330 ;
        RECT  11.960 1.745 13.765 2.125 ;
        RECT  10.465 3.090 12.325 3.330 ;
        RECT  11.960 1.100 12.325 3.330 ;
        RECT  10.465 2.640 10.805 3.330 ;
        RECT  9.015 2.640 10.805 2.920 ;
        RECT  9.015 2.640 9.365 3.190 ;
        RECT  0.375 2.640 10.805 2.915 ;
        RECT  7.560 2.640 7.930 3.185 ;
        RECT  6.135 2.640 6.475 3.190 ;
        RECT  4.695 2.640 5.040 3.175 ;
        RECT  0.375 2.640 5.040 2.920 ;
        RECT  3.255 2.640 3.595 3.190 ;
        RECT  1.815 2.640 2.155 3.200 ;
        RECT  0.375 2.640 0.715 3.185 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.000 4.100 ;
        RECT  12.705 2.630 13.045 4.100 ;
        RECT  11.225 3.560 11.565 4.100 ;
        RECT  9.745 3.165 10.085 4.100 ;
        RECT  8.295 3.150 8.635 4.100 ;
        RECT  6.855 3.145 7.195 4.100 ;
        RECT  5.415 3.150 5.755 4.100 ;
        RECT  3.975 3.150 4.315 4.100 ;
        RECT  2.535 3.150 2.875 4.100 ;
        RECT  1.095 3.150 1.435 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.000 0.180 ;
        RECT  3.255 -0.180 3.595 0.970 ;
        RECT  1.815 -0.180 2.155 0.970 ;
        RECT  0.375 -0.180 0.715 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.975 0.630 7.210 0.925 ;
        RECT  1.095 0.685 1.435 1.440 ;
        RECT  2.535 0.685 2.875 1.440 ;
        RECT  3.975 0.630 4.315 1.440 ;
        RECT  1.095 1.200 4.315 1.440 ;
        RECT  4.695 1.155 10.805 1.435 ;
        RECT  8.285 0.630 12.965 0.870 ;
        RECT  8.285 0.630 11.525 0.925 ;
        RECT  11.185 0.630 11.525 1.385 ;
        RECT  12.625 0.630 12.965 1.385 ;
    END
END NAND4T_X6_18_SVT_WB

MACRO NAND4T_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.940 1.615 8.265 2.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.360 2.320 6.710 2.660 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.080 2.320 4.500 2.660 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.105  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.995 2.320 2.460 2.695 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.129  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.080 2.945 8.820 3.285 ;
        RECT  8.495 1.045 8.820 3.285 ;
        RECT  7.720 1.045 8.820 1.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  4.800 3.515 5.140 4.100 ;
        RECT  1.840 3.515 2.180 4.100 ;
        RECT  0.370 3.125 0.670 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  1.840 -0.180 2.180 0.875 ;
        RECT  0.355 -0.180 0.690 1.020 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.600 0.520 4.400 0.815 ;
        RECT  1.080 0.535 1.420 1.345 ;
        RECT  2.600 0.520 2.940 1.345 ;
        RECT  1.080 1.105 2.940 1.345 ;
        RECT  3.320 1.045 6.620 1.340 ;
        RECT  5.520 0.475 8.780 0.815 ;
        RECT  7.000 0.475 7.340 1.340 ;
    END
END NAND4T_X4_18_SVT_WB

MACRO NAND4T_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.560 1.620 4.900 2.470 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.585  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.695 2.375 4.165 2.705 ;
        RECT  3.825 1.840 4.165 2.705 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.585  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.155 1.200 3.495 1.960 ;
        RECT  1.125 1.200 3.495 1.540 ;
        RECT  1.125 1.200 1.465 2.035 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.585  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.695 1.770 2.235 2.145 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.746  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.545 2.940 5.360 3.280 ;
        RECT  5.130 0.580 5.360 3.280 ;
        RECT  4.785 0.580 5.360 1.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.825 3.515 5.165 4.100 ;
        RECT  3.305 3.515 3.645 4.100 ;
        RECT  1.825 3.125 2.165 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  2.075 -0.180 2.415 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.215 0.580 4.405 0.920 ;
    END
END NAND4T_X2_18_SVT_WB

MACRO NAND4T_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.292  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.620 2.150 2.280 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.210 2.910 1.960 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.292  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.040 2.305 1.540 2.710 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.292  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.873  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.940 3.480 3.280 ;
        RECT  3.140 1.100 3.480 3.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.180 3.515 3.520 4.100 ;
        RECT  1.660 3.510 2.000 4.100 ;
        RECT  0.180 2.890 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.180 -0.180 0.520 1.440 ;
        END
    END VSS
END NAND4T_X1_18_SVT_WB

MACRO NAND4T_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 36.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  30.540 1.810 34.000 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.002  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  20.390 2.265 29.355 2.660 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.148  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.335 2.265 19.420 2.660 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.075  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.030 2.265 10.105 2.660 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 12.753  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  30.070 2.380 34.730 2.720 ;
        RECT  34.390 0.995 34.730 2.720 ;
        RECT  30.070 0.995 34.730 1.335 ;
        RECT  0.550 2.890 30.410 3.230 ;
        RECT  30.070 2.380 30.410 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 36.400 4.100 ;
        RECT  35.110 3.110 35.450 4.100 ;
        RECT  33.670 3.110 34.010 4.100 ;
        RECT  32.230 3.125 32.570 4.100 ;
        RECT  30.790 3.125 31.130 4.100 ;
        RECT  29.310 3.515 29.650 4.100 ;
        RECT  27.745 3.510 28.085 4.100 ;
        RECT  26.225 3.510 26.565 4.100 ;
        RECT  24.805 3.510 25.145 4.100 ;
        RECT  23.380 3.510 23.720 4.100 ;
        RECT  21.790 3.510 22.130 4.100 ;
        RECT  20.335 3.510 20.675 4.100 ;
        RECT  19.150 3.515 19.490 4.100 ;
        RECT  17.265 3.510 17.605 4.100 ;
        RECT  15.870 3.510 16.210 4.100 ;
        RECT  14.445 3.510 14.785 4.100 ;
        RECT  13.310 3.515 13.650 4.100 ;
        RECT  10.350 3.515 10.690 4.100 ;
        RECT  8.830 3.515 9.170 4.100 ;
        RECT  7.310 3.460 7.650 4.100 ;
        RECT  5.790 3.515 6.130 4.100 ;
        RECT  4.270 3.515 4.610 4.100 ;
        RECT  1.310 3.515 1.650 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 36.400 0.180 ;
        RECT  9.590 -0.180 9.930 0.795 ;
        RECT  8.070 -0.180 8.410 0.810 ;
        RECT  6.550 -0.180 6.890 0.810 ;
        RECT  5.030 -0.180 5.370 0.810 ;
        RECT  3.510 -0.180 3.850 0.810 ;
        RECT  2.070 -0.180 2.410 0.810 ;
        RECT  0.550 -0.180 0.890 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.270 1.100 1.610 1.845 ;
        RECT  1.270 1.505 19.530 1.845 ;
        RECT  11.110 0.470 20.250 0.810 ;
        RECT  19.910 0.470 20.250 1.280 ;
        RECT  19.910 0.995 28.890 1.280 ;
        RECT  20.630 0.470 35.530 0.765 ;
    END
END NAND4T_X16_18_SVT_WB

MACRO NAND4T_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.355 1.805 18.885 2.145 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.626  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.365 2.265 16.470 2.660 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.772  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.185 2.265 11.085 2.660 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.699  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.885 2.265 5.445 2.660 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.945  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.885 2.380 20.105 2.720 ;
        RECT  19.765 1.040 20.105 2.720 ;
        RECT  16.885 1.040 20.105 1.380 ;
        RECT  0.405 2.890 17.225 3.230 ;
        RECT  16.885 2.380 17.225 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 21.280 4.100 ;
        RECT  20.485 3.110 20.825 4.100 ;
        RECT  19.045 3.110 19.385 4.100 ;
        RECT  17.605 3.125 17.945 4.100 ;
        RECT  16.125 3.515 16.465 4.100 ;
        RECT  14.605 3.515 14.945 4.100 ;
        RECT  13.085 3.515 13.425 4.100 ;
        RECT  10.125 3.515 10.465 4.100 ;
        RECT  8.605 3.515 8.945 4.100 ;
        RECT  5.645 3.515 5.985 4.100 ;
        RECT  4.125 3.515 4.465 4.100 ;
        RECT  1.165 3.515 1.505 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 21.280 0.180 ;
        RECT  4.885 -0.180 5.225 0.810 ;
        RECT  3.365 -0.180 3.705 0.810 ;
        RECT  1.925 -0.180 2.265 0.810 ;
        RECT  0.405 -0.180 0.745 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.125 1.100 1.465 1.845 ;
        RECT  1.125 1.505 10.425 1.845 ;
        RECT  6.405 0.470 11.225 0.810 ;
        RECT  10.885 0.470 11.225 1.380 ;
        RECT  10.885 1.040 15.705 1.380 ;
        RECT  11.605 0.470 20.825 0.810 ;
    END
END NAND4T_X12_18_SVT_WB

MACRO NAND4T_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND4T_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.565 2.785 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.330 2.320 2.660 ;
        RECT  1.770 2.330 2.040 2.850 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.260 1.650 1.870 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.690 0.980 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.015 1.010 3.245 3.270 ;
        RECT  2.270 2.890 3.245 3.270 ;
        RECT  2.820 1.010 3.245 1.335 ;
        RECT  0.900 3.080 2.560 3.420 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 3.080 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.400 -0.180 0.740 0.930 ;
        END
    END VSS
END NAND4T_X0_18_SVT_WB

MACRO NAND3_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.290 1.820 8.100 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.170 1.360 5.510 1.950 ;
        RECT  0.700 1.360 5.510 1.590 ;
        RECT  2.660 1.360 3.470 1.905 ;
        RECT  0.700 1.360 3.470 1.630 ;
        RECT  0.700 1.360 1.060 2.150 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.420 2.135 4.700 2.365 ;
        RECT  3.890 1.820 4.700 2.365 ;
        RECT  1.420 1.860 2.230 2.365 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.860  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.720 2.695 8.060 3.395 ;
        RECT  6.080 1.105 7.860 1.440 ;
        RECT  6.370 2.695 8.060 3.035 ;
        RECT  6.370 1.105 6.710 3.395 ;
        RECT  5.210 2.180 6.710 2.410 ;
        RECT  6.080 1.105 6.710 1.540 ;
        RECT  4.930 2.695 5.440 3.395 ;
        RECT  5.210 2.180 5.440 3.395 ;
        RECT  0.940 2.695 5.440 2.925 ;
        RECT  3.610 2.695 3.950 3.395 ;
        RECT  2.280 2.695 2.620 3.395 ;
        RECT  0.940 2.695 1.280 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.440 2.655 8.780 4.100 ;
        RECT  5.670 2.640 5.990 4.100 ;
        RECT  0.220 2.475 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  4.170 -0.180 4.510 0.360 ;
        RECT  1.700 -0.180 2.040 0.360 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.500 0.535 0.840 0.875 ;
        RECT  0.500 0.590 8.580 0.875 ;
        RECT  8.240 0.590 8.580 1.345 ;
    END
END NAND3_X8_18_SVT_WB

MACRO NAND3_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.450 1.615 6.060 2.290 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.135 4.340 2.365 ;
        RECT  3.770 1.770 4.340 2.365 ;
        RECT  1.750 1.915 2.090 2.365 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.990 1.455 3.330 1.905 ;
        RECT  0.660 1.455 3.330 1.685 ;
        RECT  0.660 1.455 1.000 2.305 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.107  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 2.625 6.540 3.380 ;
        RECT  4.620 1.100 6.540 1.385 ;
        RECT  6.200 0.630 6.540 1.385 ;
        RECT  0.900 2.625 6.540 3.020 ;
        RECT  4.880 2.625 5.220 3.380 ;
        RECT  4.620 1.100 4.900 3.020 ;
        RECT  3.550 2.625 3.890 3.380 ;
        RECT  2.230 2.625 2.570 3.380 ;
        RECT  0.900 2.625 1.240 3.380 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  0.180 2.680 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  2.770 -0.180 3.110 0.740 ;
        RECT  0.180 -0.180 0.520 1.225 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.860 0.575 5.760 0.870 ;
        RECT  3.860 0.575 4.200 1.225 ;
        RECT  1.620 0.970 4.200 1.225 ;
    END
END NAND3_X6_18_SVT_WB

MACRO NAND3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.635 2.660 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.360 1.095 3.700 1.980 ;
        RECT  1.260 1.095 3.700 1.405 ;
        RECT  1.260 1.095 1.620 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.610 2.380 4.370 2.720 ;
        RECT  4.030 1.860 4.370 2.720 ;
        RECT  0.610 1.840 0.950 2.720 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.760 3.045 4.915 3.295 ;
        RECT  4.600 0.635 4.915 3.295 ;
        RECT  2.320 0.635 4.915 0.865 ;
        RECT  2.320 0.470 2.660 0.865 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.080 3.560 3.420 4.100 ;
        RECT  1.560 3.560 1.900 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.520 -0.180 4.860 0.405 ;
        RECT  0.180 -0.180 0.520 1.280 ;
        END
    END VSS
END NAND3_X4_18_SVT_WB

MACRO NAND3_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.225 1.355 2.160 1.640 ;
        RECT  1.225 1.165 1.555 1.640 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.870 3.325 2.100 ;
        RECT  2.800 1.545 3.325 2.100 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.330 3.885 2.560 ;
        RECT  3.635 2.040 3.885 2.560 ;
        RECT  0.130 2.085 0.820 2.560 ;
        RECT  0.130 1.665 0.450 2.560 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.817  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.790 4.365 3.130 ;
        RECT  4.115 0.785 4.365 3.130 ;
        RECT  4.045 0.785 4.365 1.665 ;
        RECT  2.110 0.785 4.365 1.125 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  1.590 3.515 2.870 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.920 -0.180 4.260 0.460 ;
        RECT  0.240 -0.180 0.580 1.010 ;
        END
    END VSS
END NAND3_X3_18_SVT_WB

MACRO NAND3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.860 2.105 2.875 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.770 1.540 2.275 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.260 1.030 1.560 ;
        RECT  0.420 1.260 0.760 1.960 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.677  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 3.110 2.660 3.450 ;
        RECT  2.335 0.550 2.660 3.450 ;
        RECT  2.260 0.550 2.660 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.640 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
END NAND3_X2_18_SVT_WB

MACRO NAND3_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.960  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.810 1.615 21.825 2.135 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.960  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.090 1.040 14.440 1.995 ;
        RECT  0.655 1.040 14.440 1.270 ;
        RECT  11.450 1.040 11.820 1.905 ;
        RECT  8.570 1.040 8.930 1.905 ;
        RECT  5.690 1.040 6.060 1.905 ;
        RECT  2.805 1.040 3.180 1.905 ;
        RECT  0.655 1.040 1.010 1.910 ;
        RECT  0.655 1.040 0.945 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.960  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.120 2.135 13.095 2.365 ;
        RECT  12.525 1.630 13.095 2.365 ;
        RECT  10.000 1.640 10.565 2.365 ;
        RECT  7.050 1.640 7.610 2.365 ;
        RECT  4.240 1.705 4.625 2.365 ;
        RECT  4.315 1.655 4.545 2.365 ;
        RECT  2.120 1.670 2.510 2.365 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 12.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.290 2.435 21.400 2.665 ;
        RECT  15.010 1.155 21.110 1.385 ;
        RECT  18.055 1.155 18.410 2.665 ;
        RECT  0.900 2.705 15.640 2.935 ;
        RECT  15.290 2.435 15.640 2.935 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 22.400 4.100 ;
        RECT  21.780 3.165 22.120 4.100 ;
        RECT  20.340 3.165 20.680 4.100 ;
        RECT  18.900 3.165 19.240 4.100 ;
        RECT  17.460 3.165 17.800 4.100 ;
        RECT  16.020 3.165 16.360 4.100 ;
        RECT  14.580 3.165 14.920 4.100 ;
        RECT  13.140 3.165 13.480 4.100 ;
        RECT  11.700 3.165 12.040 4.100 ;
        RECT  10.260 3.165 10.600 4.100 ;
        RECT  8.820 3.165 9.160 4.100 ;
        RECT  7.380 3.165 7.720 4.100 ;
        RECT  5.940 3.165 6.280 4.100 ;
        RECT  4.500 3.165 4.840 4.100 ;
        RECT  3.060 3.165 3.400 4.100 ;
        RECT  1.620 3.165 1.960 4.100 ;
        RECT  0.180 3.165 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 22.400 0.180 ;
        RECT  13.100 -0.180 13.440 0.350 ;
        RECT  10.210 -0.180 10.550 0.350 ;
        RECT  7.325 -0.180 7.665 0.350 ;
        RECT  4.440 -0.180 4.780 0.350 ;
        RECT  1.815 -0.180 2.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 0.580 21.830 0.810 ;
    END
END NAND3_X24_18_SVT_WB

MACRO NAND3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.820 2.150 2.355 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 0.895 1.540 1.725 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.565 1.770 0.980 2.395 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.839  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.915 2.625 2.660 2.965 ;
        RECT  2.380 0.865 2.660 2.965 ;
        RECT  2.265 0.865 2.660 1.205 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  1.675 3.515 2.015 4.100 ;
        RECT  0.195 2.730 0.535 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.195 -0.180 0.535 1.100 ;
        END
    END VSS
END NAND3_X1_18_SVT_WB

MACRO NAND3_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.085 1.665 17.325 2.205 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.000 1.830 11.545 2.190 ;
        RECT  11.000 1.150 11.230 2.190 ;
        RECT  0.685 1.150 11.230 1.380 ;
        RECT  8.575 1.150 8.930 1.905 ;
        RECT  5.685 1.150 6.050 1.905 ;
        RECT  2.815 1.150 3.165 1.905 ;
        RECT  0.755 1.150 1.020 2.010 ;
        RECT  0.685 1.150 1.020 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.150 2.135 10.070 2.365 ;
        RECT  9.550 1.620 10.070 2.365 ;
        RECT  7.130 1.625 7.490 2.365 ;
        RECT  4.240 1.630 4.635 2.365 ;
        RECT  2.150 1.745 2.495 2.365 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.720  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.795 2.435 17.080 2.715 ;
        RECT  12.470 2.435 17.080 2.665 ;
        RECT  12.130 1.125 16.790 1.355 ;
        RECT  13.760 1.125 14.485 2.665 ;
        RECT  0.900 2.705 12.760 2.935 ;
        RECT  12.470 2.435 12.760 2.935 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  16.020 3.165 16.360 4.100 ;
        RECT  14.580 3.165 14.920 4.100 ;
        RECT  13.140 3.165 13.480 4.100 ;
        RECT  11.700 3.165 12.040 4.100 ;
        RECT  10.260 3.165 10.600 4.100 ;
        RECT  8.820 3.165 9.160 4.100 ;
        RECT  7.380 3.165 7.720 4.100 ;
        RECT  5.940 3.165 6.280 4.100 ;
        RECT  4.500 3.165 4.840 4.100 ;
        RECT  3.060 3.165 3.400 4.100 ;
        RECT  1.620 3.165 1.960 4.100 ;
        RECT  0.180 2.635 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  10.010 -0.180 10.350 0.350 ;
        RECT  7.630 -0.180 7.970 0.350 ;
        RECT  4.400 -0.180 4.755 0.350 ;
        RECT  1.800 -0.180 2.155 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.365 0.580 17.535 0.810 ;
        RECT  17.150 0.580 17.535 1.350 ;
    END
END NAND3_X16_18_SVT_WB

MACRO NAND3_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.095 1.800 12.295 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.570 1.640 8.080 1.980 ;
        RECT  7.570 1.260 7.800 1.980 ;
        RECT  2.870 1.260 7.800 1.600 ;
        RECT  5.520 1.260 5.860 1.905 ;
        RECT  2.870 1.260 5.860 1.640 ;
        RECT  2.870 1.260 3.210 1.905 ;
        RECT  0.700 1.260 7.800 1.590 ;
        RECT  0.420 1.640 0.930 1.980 ;
        RECT  0.700 1.260 0.930 1.980 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.135 7.020 2.365 ;
        RECT  6.680 1.860 7.020 2.365 ;
        RECT  4.390 1.870 4.730 2.365 ;
        RECT  1.740 1.820 2.150 2.365 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.290  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.640 2.695 11.980 3.395 ;
        RECT  8.975 1.105 11.890 1.400 ;
        RECT  10.290 2.695 11.980 2.980 ;
        RECT  10.290 2.695 10.630 3.395 ;
        RECT  0.900 2.695 11.980 2.925 ;
        RECT  8.975 1.105 9.630 2.925 ;
        RECT  8.850 2.695 9.190 3.450 ;
        RECT  8.670 1.105 11.890 1.385 ;
        RECT  7.520 2.695 7.860 3.450 ;
        RECT  6.200 2.695 6.540 3.450 ;
        RECT  4.870 2.695 5.210 3.450 ;
        RECT  3.550 2.695 3.890 3.450 ;
        RECT  2.220 2.695 2.560 3.450 ;
        RECT  0.900 2.695 1.240 3.400 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  12.360 2.695 12.700 4.100 ;
        RECT  0.180 2.475 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  6.670 -0.180 7.010 0.360 ;
        RECT  4.110 -0.180 4.450 0.360 ;
        RECT  1.460 -0.180 1.800 0.360 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.535 0.520 0.875 ;
        RECT  0.180 0.590 12.610 0.875 ;
        RECT  12.270 0.590 12.610 1.345 ;
    END
END NAND3_X12_18_SVT_WB

MACRO NAND3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.570 2.150 2.190 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.065 1.540 1.590 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.810 1.030 2.355 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.727  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.585 2.660 2.925 ;
        RECT  2.380 0.730 2.660 2.925 ;
        RECT  2.240 0.730 2.660 1.070 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  1.660 3.515 2.000 4.100 ;
        RECT  0.180 2.585 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.230 -0.180 0.570 1.070 ;
        END
    END VSS
END NAND3_X0_18_SVT_WB

MACRO NAND3T_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.960 1.615 9.455 2.540 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.437  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.380 1.675 8.730 2.305 ;
        RECT  1.335 1.675 8.730 1.905 ;
        RECT  5.790 1.675 6.660 2.285 ;
        RECT  3.420 1.675 4.240 2.345 ;
        RECT  0.775 2.210 1.570 2.550 ;
        RECT  1.335 1.675 1.565 2.550 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.248  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.275 2.650 7.795 2.880 ;
        RECT  6.960 2.240 7.795 2.880 ;
        RECT  4.555 2.235 5.410 2.880 ;
        RECT  2.275 2.280 3.125 2.880 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.992  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.985 1.760 11.365 2.880 ;
        RECT  11.000 1.155 11.365 2.880 ;
        RECT  9.715 1.760 11.365 2.150 ;
        RECT  1.040 3.110 9.980 3.340 ;
        RECT  9.715 1.760 9.980 3.340 ;
        RECT  9.715 1.155 9.945 3.340 ;
        RECT  9.570 1.155 9.945 1.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.800 2.640 12.140 4.100 ;
        RECT  10.360 2.635 10.700 4.100 ;
        RECT  3.120 3.570 3.460 4.100 ;
        RECT  0.320 3.110 0.660 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  7.245 -0.180 7.595 0.350 ;
        RECT  4.865 -0.180 5.215 0.350 ;
        RECT  2.490 -0.180 2.830 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.275 1.040 2.100 1.270 ;
        RECT  0.990 0.580 12.070 0.810 ;
        RECT  10.275 0.580 10.645 1.280 ;
        RECT  3.660 0.580 4.030 1.285 ;
        RECT  6.040 0.580 6.410 1.285 ;
        RECT  8.740 0.580 9.130 1.335 ;
        RECT  11.740 0.580 12.070 1.335 ;
    END
END NAND3T_X8_18_SVT_WB

MACRO NAND3T_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.390 1.705 8.190 2.085 ;
        RECT  7.390 1.705 7.755 2.185 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.728  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.180 1.760 6.990 2.340 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.782  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.765 3.210 2.280 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.107  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.615 2.375 9.845 3.190 ;
        RECT  8.520 1.100 9.845 1.455 ;
        RECT  9.615 0.630 9.845 1.455 ;
        RECT  8.120 2.375 9.845 2.700 ;
        RECT  8.520 1.100 8.840 2.700 ;
        RECT  8.175 1.100 9.845 1.445 ;
        RECT  8.120 2.375 8.405 3.190 ;
        RECT  0.920 2.595 8.405 2.825 ;
        RECT  6.680 2.595 7.035 3.320 ;
        RECT  5.240 2.595 5.590 3.220 ;
        RECT  3.805 2.595 4.145 3.190 ;
        RECT  2.350 2.595 2.710 3.190 ;
        RECT  0.920 2.595 1.260 3.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  8.840 3.105 9.180 4.100 ;
        RECT  7.400 3.110 7.740 4.100 ;
        RECT  5.960 3.105 6.300 4.100 ;
        RECT  4.520 3.105 4.860 4.100 ;
        RECT  3.080 3.055 3.420 4.100 ;
        RECT  1.645 3.095 1.980 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  3.040 -0.180 3.380 0.405 ;
        RECT  1.515 -0.180 1.865 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.760 0.635 7.020 0.865 ;
        RECT  3.805 0.635 4.140 1.400 ;
        RECT  2.260 0.635 2.630 1.420 ;
        RECT  0.760 0.635 1.105 1.425 ;
        RECT  7.455 0.515 9.180 0.755 ;
        RECT  7.455 0.515 7.685 1.435 ;
        RECT  4.505 1.095 7.685 1.435 ;
    END
END NAND3T_X6_18_SVT_WB

MACRO NAND3T_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.170 1.675 5.765 2.400 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.058  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.485 2.060 4.940 2.400 ;
        RECT  2.755 2.640 4.715 2.870 ;
        RECT  4.485 2.060 4.715 2.870 ;
        RECT  2.240 2.125 3.075 2.675 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.285  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.385 2.120 4.230 2.405 ;
        RECT  3.385 1.575 3.680 2.405 ;
        RECT  1.315 1.575 3.680 1.835 ;
        RECT  0.810 2.145 1.630 2.675 ;
        RECT  1.315 1.575 1.630 2.675 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.825  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.475 3.100 6.585 3.330 ;
        RECT  6.040 1.100 6.585 3.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.815 2.545 7.100 4.100 ;
        RECT  5.250 3.560 5.590 4.100 ;
        RECT  0.730 2.955 1.090 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  3.635 -0.180 3.975 0.885 ;
        RECT  1.045 -0.180 1.385 0.790 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.325 0.470 0.655 1.250 ;
        RECT  0.325 1.020 2.120 1.250 ;
        RECT  5.125 0.630 7.100 0.870 ;
        RECT  5.125 0.630 5.490 1.345 ;
        RECT  2.455 1.115 5.490 1.345 ;
        RECT  6.815 0.630 7.100 1.440 ;
    END
END NAND3T_X4_18_SVT_WB

MACRO NAND3T_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.960 1.735 4.340 2.270 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.585  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.765 1.770 3.700 2.270 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.585  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.555 2.000 2.200 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.600 2.500 4.900 2.840 ;
        RECT  4.570 0.630 4.900 2.840 ;
        RECT  4.280 2.500 4.620 3.200 ;
        RECT  2.600 2.500 2.940 3.255 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.520 3.070 3.860 4.100 ;
        RECT  1.740 2.555 2.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.660 -0.180 2.000 0.400 ;
        RECT  0.180 -0.180 0.520 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.630 3.445 0.920 ;
        RECT  0.900 0.535 1.240 1.325 ;
        RECT  3.800 0.685 4.140 1.440 ;
        RECT  2.330 1.150 4.140 1.440 ;
    END
END NAND3T_X2_18_SVT_WB

MACRO NAND3T_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.090 2.100 1.625 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.292  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.340 1.650 2.775 ;
        RECT  1.210 1.965 1.520 2.775 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.292  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.620 0.980 2.430 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.839  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.940 3.110 2.660 3.450 ;
        RECT  2.330 0.520 2.660 3.450 ;
        RECT  1.970 0.520 2.660 0.860 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.955 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.220 -0.180 0.560 1.330 ;
        END
    END VSS
END NAND3T_X1_18_SVT_WB

MACRO NAND3T_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.865 1.820 23.375 2.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.412  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  18.285 1.820 18.630 2.160 ;
        RECT  2.015 1.820 18.630 2.090 ;
        RECT  15.685 1.820 16.495 2.180 ;
        RECT  13.275 1.820 13.615 2.180 ;
        RECT  10.565 1.820 11.375 2.180 ;
        RECT  7.605 1.820 8.415 2.180 ;
        RECT  4.870 1.820 5.680 2.180 ;
        RECT  2.015 1.820 2.825 2.180 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.847  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.410 17.670 2.660 ;
        RECT  16.860 2.320 17.670 2.660 ;
        RECT  14.460 2.320 15.300 2.660 ;
        RECT  12.000 2.320 12.810 2.660 ;
        RECT  9.130 2.320 9.940 2.660 ;
        RECT  6.185 2.320 6.995 2.660 ;
        RECT  3.535 2.320 4.345 2.660 ;
        RECT  0.650 2.320 1.470 2.660 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.818  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  23.605 1.145 24.180 2.935 ;
        RECT  19.425 2.595 24.180 2.935 ;
        RECT  19.230 1.145 24.180 1.440 ;
        RECT  0.900 2.890 19.860 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 25.200 4.100 ;
        RECT  24.560 3.065 24.900 4.100 ;
        RECT  23.120 3.165 23.460 4.100 ;
        RECT  21.680 3.165 22.020 4.100 ;
        RECT  20.240 3.165 20.580 4.100 ;
        RECT  13.000 3.510 13.340 4.100 ;
        RECT  8.600 3.510 8.940 4.100 ;
        RECT  3.005 3.510 3.345 4.100 ;
        RECT  0.180 3.105 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 25.200 0.180 ;
        RECT  17.140 -0.180 17.480 0.405 ;
        RECT  14.685 -0.180 15.025 0.405 ;
        RECT  12.280 -0.180 12.620 0.405 ;
        RECT  6.465 -0.180 6.805 0.405 ;
        RECT  3.805 -0.180 4.145 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 0.520 1.545 ;
        RECT  0.180 1.205 3.305 1.545 ;
        RECT  2.245 0.635 24.900 0.915 ;
        RECT  2.245 0.635 18.850 0.975 ;
        RECT  18.510 0.635 18.850 1.440 ;
        RECT  24.560 0.635 24.900 1.440 ;
        RECT  5.105 0.635 5.445 1.590 ;
        RECT  7.840 0.635 8.180 1.590 ;
        RECT  10.800 0.635 11.140 1.590 ;
        RECT  13.495 0.635 13.835 1.590 ;
        RECT  15.920 0.635 16.260 1.590 ;
    END
END NAND3T_X16_18_SVT_WB

MACRO NAND3T_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.440 1.760 15.720 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.368  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.720 1.820 14.060 2.320 ;
        RECT  0.420 1.820 14.060 2.090 ;
        RECT  11.000 1.820 11.820 2.200 ;
        RECT  8.600 1.820 8.990 2.200 ;
        RECT  5.880 1.820 6.690 2.200 ;
        RECT  3.400 1.820 3.740 2.200 ;
        RECT  0.420 1.820 0.760 2.160 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.537  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.190 2.430 12.990 2.660 ;
        RECT  12.180 2.320 12.990 2.660 ;
        RECT  9.830 2.320 10.640 2.660 ;
        RECT  7.330 2.320 8.140 2.660 ;
        RECT  4.450 2.320 5.260 2.660 ;
        RECT  2.190 2.320 2.530 2.660 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.501  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  17.800 1.145 18.140 2.935 ;
        RECT  14.920 2.640 18.140 2.935 ;
        RECT  14.910 1.145 18.140 1.440 ;
        RECT  0.200 2.895 15.260 3.235 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 19.040 4.100 ;
        RECT  18.520 2.380 18.860 4.100 ;
        RECT  17.080 3.165 17.420 4.100 ;
        RECT  15.640 3.165 15.980 4.100 ;
        RECT  12.720 3.510 13.060 4.100 ;
        RECT  8.320 3.510 8.660 4.100 ;
        RECT  3.920 3.510 4.260 4.100 ;
        RECT  0.960 3.515 1.430 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 19.040 0.180 ;
        RECT  12.540 -0.180 12.880 0.405 ;
        RECT  10.020 -0.180 10.360 0.405 ;
        RECT  7.600 -0.180 7.940 0.405 ;
        RECT  4.930 -0.180 5.270 0.405 ;
        RECT  1.970 -0.180 2.310 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 0.635 18.860 0.915 ;
        RECT  0.200 0.635 14.300 0.975 ;
        RECT  0.200 0.635 0.540 1.440 ;
        RECT  13.960 0.635 14.300 1.440 ;
        RECT  18.520 0.635 18.860 1.440 ;
        RECT  3.160 0.635 3.500 1.445 ;
        RECT  6.120 0.635 6.460 1.445 ;
        RECT  8.830 0.635 9.170 1.445 ;
        RECT  11.240 0.635 11.580 1.445 ;
    END
END NAND3T_X12_18_SVT_WB

MACRO NAND3T_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND3T_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.340 2.150 2.150 ;
        RECT  1.670 1.340 2.150 1.680 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 2.055 1.565 2.815 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.620 0.800 2.430 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.940 3.045 2.660 3.385 ;
        RECT  2.380 0.680 2.660 3.385 ;
        RECT  2.090 0.680 2.660 1.020 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 3.045 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.220 -0.180 0.560 1.020 ;
        END
    END VSS
END NAND3T_X0_18_SVT_WB

MACRO NAND2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.350 1.820 4.440 2.160 ;
        RECT  1.660 2.135 3.690 2.365 ;
        RECT  1.660 1.860 2.000 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.280 1.360 5.585 1.960 ;
        RECT  0.870 1.360 5.585 1.590 ;
        RECT  2.660 1.360 3.000 1.905 ;
        RECT  0.870 1.360 3.000 1.630 ;
        RECT  0.520 1.805 1.100 2.145 ;
        RECT  0.870 1.360 1.100 2.145 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.618  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.595 6.045 2.825 ;
        RECT  5.815 0.640 6.045 2.825 ;
        RECT  1.460 0.640 6.045 0.980 ;
        RECT  5.045 2.595 5.400 3.405 ;
        RECT  3.620 2.595 3.960 3.405 ;
        RECT  2.180 2.595 3.960 2.835 ;
        RECT  2.180 2.595 2.520 3.405 ;
        RECT  0.740 2.595 1.075 3.445 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.340 3.065 4.680 4.100 ;
        RECT  2.900 3.065 3.240 4.100 ;
        RECT  1.460 3.065 1.800 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  5.640 -0.180 5.980 0.410 ;
        RECT  2.860 -0.180 3.200 0.405 ;
        RECT  0.180 -0.180 0.520 1.440 ;
        END
    END VSS
END NAND2_X8_18_SVT_WB

MACRO NAND2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.435 1.820 4.300 2.200 ;
        RECT  1.905 2.135 3.775 2.365 ;
        RECT  1.905 1.915 2.245 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.455 3.205 1.905 ;
        RECT  0.985 1.455 3.205 1.685 ;
        RECT  0.650 1.810 1.225 2.150 ;
        RECT  0.985 1.455 1.225 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.825 2.595 4.825 2.935 ;
        RECT  4.535 0.630 4.825 2.935 ;
        RECT  4.530 0.995 4.825 2.935 ;
        RECT  1.665 0.995 4.825 1.225 ;
        RECT  3.825 2.595 4.165 3.405 ;
        RECT  0.945 2.595 4.825 2.835 ;
        RECT  2.380 2.595 2.725 3.405 ;
        RECT  0.945 2.595 2.725 2.935 ;
        RECT  1.665 0.885 2.005 1.225 ;
        RECT  0.945 2.595 1.285 3.410 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.105 3.065 3.445 4.100 ;
        RECT  1.665 3.165 2.005 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.105 -0.180 3.445 0.765 ;
        RECT  0.225 -0.180 0.565 1.280 ;
        END
    END VSS
END NAND2_X6_18_SVT_WB

MACRO NAND2_X5_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.988  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.880 2.155 4.390 2.395 ;
        RECT  4.010 1.820 4.390 2.395 ;
        RECT  1.880 2.055 2.220 2.395 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.988  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.600 1.595 2.940 1.925 ;
        RECT  0.650 1.595 2.940 1.825 ;
        RECT  0.650 1.595 1.030 2.100 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.440  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.920 2.640 4.860 2.880 ;
        RECT  4.620 1.025 4.860 2.880 ;
        RECT  1.640 1.135 4.860 1.365 ;
        RECT  4.520 1.025 4.860 1.365 ;
        RECT  3.800 2.640 4.140 3.450 ;
        RECT  2.360 2.640 2.700 3.450 ;
        RECT  1.640 1.025 1.980 1.365 ;
        RECT  0.920 2.640 1.260 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.520 3.110 4.860 4.100 ;
        RECT  3.080 3.110 3.420 4.100 ;
        RECT  1.640 3.110 1.980 4.100 ;
        RECT  0.200 2.640 0.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.080 -0.180 3.420 0.905 ;
        RECT  0.450 -0.180 0.790 1.345 ;
        END
    END VSS
END NAND2_X5_18_SVT_WB

MACRO NAND2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.635 2.150 2.140 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.550 2.370 2.785 2.710 ;
        RECT  2.450 1.860 2.785 2.710 ;
        RECT  0.550 1.860 0.890 2.710 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.893  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.940 3.245 3.330 ;
        RECT  3.015 1.065 3.245 3.330 ;
        RECT  1.540 1.065 3.245 1.405 ;
        RECT  1.540 0.595 1.880 1.405 ;
        RECT  0.740 2.940 1.080 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.500 3.560 1.840 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.690 -0.180 3.030 0.810 ;
        RECT  0.310 -0.180 0.650 1.290 ;
        END
    END VSS
END NAND2_X4_18_SVT_WB

MACRO NAND2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.210 1.745 1.695 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.685 1.925 2.775 2.165 ;
        RECT  2.435 1.825 2.775 2.165 ;
        RECT  0.685 1.770 1.025 2.165 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.353  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.925 2.820 3.245 3.160 ;
        RECT  3.005 0.640 3.245 3.160 ;
        RECT  1.525 0.640 3.245 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 2.380 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.205 -0.180 0.545 1.175 ;
        END
    END VSS
END NAND2_X3_18_SVT_WB

MACRO NAND2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.175 1.595 1.540 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.460 2.335 1.030 2.675 ;
        RECT  0.460 1.840 0.850 2.675 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.940 2.905 2.100 3.245 ;
        RECT  1.770 0.470 2.100 3.245 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.700 3.475 2.040 4.100 ;
        RECT  0.220 3.125 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.180 -0.180 0.520 1.440 ;
        END
    END VSS
END NAND2_X2_18_SVT_WB

MACRO NAND2_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.752  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.580 2.135 15.670 2.365 ;
        RECT  15.280 1.820 15.670 2.365 ;
        RECT  12.450 1.860 12.790 2.365 ;
        RECT  10.050 1.860 10.390 2.365 ;
        RECT  6.810 1.820 7.200 2.365 ;
        RECT  3.980 1.860 4.320 2.365 ;
        RECT  1.580 1.860 1.920 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.752  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.480 1.360 16.765 2.185 ;
        RECT  9.230 1.360 16.765 1.590 ;
        RECT  13.650 1.360 13.990 1.905 ;
        RECT  9.230 1.360 13.990 1.630 ;
        RECT  11.490 1.360 11.830 1.905 ;
        RECT  8.005 1.620 9.570 1.905 ;
        RECT  8.005 1.210 8.380 1.905 ;
        RECT  0.760 1.360 8.380 1.590 ;
        RECT  7.980 1.210 8.380 1.590 ;
        RECT  5.180 1.360 5.520 1.905 ;
        RECT  0.760 1.360 5.520 1.630 ;
        RECT  3.020 1.360 3.360 1.905 ;
        RECT  0.260 1.620 1.100 1.960 ;
        RECT  0.260 1.620 0.545 2.010 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 10.860  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.640 17.245 2.880 ;
        RECT  16.995 0.635 17.245 2.880 ;
        RECT  1.320 0.635 17.245 0.980 ;
        RECT  16.175 2.640 16.535 3.450 ;
        RECT  14.850 2.640 15.190 3.450 ;
        RECT  13.410 2.640 13.750 3.450 ;
        RECT  11.970 2.640 12.310 3.450 ;
        RECT  10.530 2.640 10.870 3.450 ;
        RECT  9.210 2.640 9.550 3.420 ;
        RECT  7.820 2.640 8.160 3.450 ;
        RECT  6.380 2.640 6.720 3.450 ;
        RECT  4.940 2.640 5.280 3.450 ;
        RECT  3.500 2.640 3.840 3.450 ;
        RECT  2.060 2.640 2.400 3.450 ;
        RECT  0.740 2.640 1.080 3.420 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.360 4.100 ;
        RECT  14.130 3.110 14.470 4.100 ;
        RECT  12.690 3.110 13.030 4.100 ;
        RECT  11.250 3.110 11.590 4.100 ;
        RECT  7.100 3.110 7.440 4.100 ;
        RECT  5.660 3.110 6.000 4.100 ;
        RECT  4.220 3.110 4.560 4.100 ;
        RECT  2.780 3.110 3.120 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.360 0.180 ;
        RECT  16.760 -0.180 17.100 0.405 ;
        RECT  14.090 -0.180 14.430 0.405 ;
        RECT  11.290 -0.180 11.630 0.405 ;
        RECT  8.290 -0.180 8.635 0.405 ;
        RECT  5.620 -0.180 5.960 0.405 ;
        RECT  2.820 -0.180 3.160 0.405 ;
        RECT  0.190 -0.180 0.530 1.390 ;
        END
    END VSS
END NAND2_X24_18_SVT_WB

MACRO NAND2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.310 1.175 1.540 1.660 ;
        RECT  1.090 1.175 1.540 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.525 1.820 1.030 2.135 ;
        RECT  0.525 1.685 0.860 2.135 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.562  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.000 2.380 2.100 2.660 ;
        RECT  1.770 0.605 2.100 2.660 ;
        RECT  1.705 0.605 2.100 0.945 ;
        RECT  1.000 2.380 1.340 3.020 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.720 2.890 2.060 4.100 ;
        RECT  0.280 2.680 0.620 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.280 -0.180 0.620 1.050 ;
        END
    END VSS
END NAND2_X1_18_SVT_WB

MACRO NAND2_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.710 1.865 9.995 2.145 ;
        RECT  9.430 1.915 9.995 2.145 ;
        RECT  2.760 2.135 9.660 2.365 ;
        RECT  6.940 1.915 7.280 2.365 ;
        RECT  3.980 1.915 4.320 2.365 ;
        RECT  2.760 1.820 2.990 2.365 ;
        RECT  1.620 1.820 2.990 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.225 1.615 11.135 1.965 ;
        RECT  10.225 1.360 10.455 1.965 ;
        RECT  0.930 1.360 10.455 1.590 ;
        RECT  8.090 1.360 8.430 1.905 ;
        RECT  5.420 1.360 5.760 1.905 ;
        RECT  3.310 1.360 3.650 1.905 ;
        RECT  0.460 1.625 1.160 2.100 ;
        RECT  0.930 1.360 1.160 2.100 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.715 2.595 11.620 2.830 ;
        RECT  11.365 0.790 11.620 2.830 ;
        RECT  11.240 2.195 11.620 2.830 ;
        RECT  1.460 0.790 11.620 1.020 ;
        RECT  10.715 2.595 10.945 3.360 ;
        RECT  0.740 2.595 11.620 2.825 ;
        RECT  9.395 2.595 9.625 3.405 ;
        RECT  7.955 2.595 8.185 3.405 ;
        RECT  6.515 2.595 6.745 3.405 ;
        RECT  4.995 2.595 5.225 3.405 ;
        RECT  3.555 2.595 3.785 3.405 ;
        RECT  2.115 2.595 2.345 3.360 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  8.620 3.110 8.960 4.100 ;
        RECT  7.180 3.110 7.520 4.100 ;
        RECT  5.660 3.110 6.080 4.100 ;
        RECT  4.220 3.110 4.560 4.100 ;
        RECT  2.780 3.110 3.120 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  11.120 -0.180 11.475 0.405 ;
        RECT  8.575 -0.180 8.925 0.405 ;
        RECT  5.695 -0.180 6.040 0.405 ;
        RECT  2.815 -0.180 3.170 0.405 ;
        RECT  0.215 -0.180 0.560 1.280 ;
        END
    END VSS
END NAND2_X16_18_SVT_WB

MACRO NAND2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.580 2.135 7.200 2.365 ;
        RECT  6.810 1.820 7.200 2.365 ;
        RECT  3.980 1.860 4.320 2.365 ;
        RECT  1.580 1.860 1.920 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.040 1.205 8.380 2.185 ;
        RECT  0.760 1.360 8.380 1.590 ;
        RECT  7.980 1.205 8.380 1.590 ;
        RECT  5.180 1.360 5.520 1.905 ;
        RECT  0.760 1.360 5.520 1.630 ;
        RECT  3.020 1.360 3.360 1.905 ;
        RECT  0.260 1.620 1.100 1.960 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.640 8.845 2.870 ;
        RECT  8.610 0.635 8.845 2.870 ;
        RECT  1.340 0.635 8.845 0.975 ;
        RECT  7.820 2.640 8.160 3.450 ;
        RECT  0.740 2.640 8.160 2.880 ;
        RECT  6.380 2.640 6.720 3.450 ;
        RECT  4.940 2.640 5.280 3.450 ;
        RECT  3.500 2.640 3.840 3.450 ;
        RECT  2.060 2.640 2.400 3.450 ;
        RECT  0.740 2.640 2.400 2.980 ;
        RECT  0.740 2.640 1.080 3.420 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  7.100 3.110 7.440 4.100 ;
        RECT  5.660 3.110 6.000 4.100 ;
        RECT  4.220 3.110 4.560 4.100 ;
        RECT  2.780 3.110 3.120 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.290 -0.180 8.630 0.405 ;
        RECT  5.620 -0.180 5.960 0.405 ;
        RECT  2.820 -0.180 3.160 0.405 ;
        RECT  0.190 -0.180 0.530 1.390 ;
        END
    END VSS
END NAND2_X12_18_SVT_WB

MACRO NAND2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.120 1.070 1.540 1.605 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.820 1.030 2.100 ;
        RECT  0.520 1.540 0.860 2.100 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.000 2.330 2.105 2.670 ;
        RECT  1.770 0.510 2.105 2.670 ;
        RECT  1.660 0.510 2.105 0.840 ;
        RECT  1.000 2.330 1.340 3.240 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.720 2.900 2.060 4.100 ;
        RECT  0.280 2.900 0.620 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.280 -0.180 0.620 0.850 ;
        END
    END VSS
END NAND2_X0_18_SVT_WB

MACRO NAND2_A_OAI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_OAI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.197  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.665 0.700 2.090 ;
        RECT  0.130 1.665 0.420 2.320 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.197  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.930 1.900 1.565 2.710 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.355 1.670 2.810 2.380 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.620 3.830 2.235 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.268  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.680 2.500 8.020 3.245 ;
        RECT  7.180 0.655 8.020 1.355 ;
        RECT  6.160 2.540 8.020 2.840 ;
        RECT  7.180 2.500 8.020 2.840 ;
        RECT  7.180 0.655 7.560 2.840 ;
        RECT  6.160 0.655 8.020 1.225 ;
        RECT  6.160 2.540 6.500 3.300 ;
        RECT  6.160 0.470 6.500 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.400 2.545 8.795 4.100 ;
        RECT  6.920 3.070 7.260 4.100 ;
        RECT  5.400 3.510 5.740 4.100 ;
        RECT  3.790 3.515 4.130 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.400 -0.180 8.795 1.355 ;
        RECT  6.920 -0.180 7.260 0.410 ;
        RECT  5.400 -0.180 5.740 0.405 ;
        RECT  0.790 -0.180 1.600 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 1.105 1.425 1.435 ;
        RECT  1.085 1.105 1.425 1.670 ;
        RECT  1.085 1.440 2.080 1.670 ;
        RECT  1.795 1.440 2.080 3.385 ;
        RECT  0.870 3.045 2.080 3.385 ;
        RECT  1.995 0.530 3.800 0.870 ;
        RECT  2.740 1.100 3.270 1.440 ;
        RECT  4.380 1.840 4.885 2.180 ;
        RECT  3.040 1.100 3.270 2.950 ;
        RECT  3.040 2.575 4.610 2.950 ;
        RECT  4.380 1.840 4.610 2.950 ;
        RECT  2.310 2.610 4.610 2.950 ;
        RECT  2.310 2.610 2.650 3.385 ;
        RECT  4.840 1.100 5.345 1.440 ;
        RECT  5.115 1.860 6.675 2.200 ;
        RECT  5.115 1.100 5.345 2.735 ;
        RECT  4.840 2.410 5.345 2.735 ;
    END
END NAND2_A_OAI21_X8_18_SVT_WB

MACRO NAND2_A_OAI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_OAI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.650 0.990 2.150 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.685 1.555 2.290 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.455 4.950 2.100 ;
        RECT  2.860 1.455 4.950 1.685 ;
        RECT  2.860 1.455 3.145 1.960 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.915 3.900 2.660 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.658  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.180 0.995 5.460 2.720 ;
        RECT  2.400 0.995 5.460 1.225 ;
        RECT  2.400 2.380 2.865 2.720 ;
        RECT  2.400 0.995 2.630 2.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  6.150 2.490 6.490 4.100 ;
        RECT  3.720 3.510 4.060 4.100 ;
        RECT  1.765 3.515 2.105 4.100 ;
        RECT  0.255 2.435 0.595 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  5.875 -0.180 6.215 1.375 ;
        RECT  1.515 -0.180 1.855 0.955 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.275 0.470 5.495 0.765 ;
        RECT  0.255 0.670 0.595 1.420 ;
        RECT  0.255 1.190 2.170 1.420 ;
        RECT  1.885 1.190 2.170 3.180 ;
        RECT  0.975 2.840 2.170 3.180 ;
        RECT  5.690 1.840 5.920 3.180 ;
        RECT  0.975 2.950 5.920 3.180 ;
        RECT  0.975 2.575 1.315 3.385 ;
    END
END NAND2_A_OAI21_X4_18_SVT_WB

MACRO NAND2_A_OAI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_OAI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.630 0.600 2.275 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.050 2.290 1.540 2.710 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.125 2.725 2.395 ;
        RECT  2.380 1.770 2.725 2.395 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.770 3.780 2.450 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.680 1.100 3.300 1.540 ;
        RECT  2.265 2.640 3.185 2.935 ;
        RECT  2.955 1.100 3.185 2.935 ;
        RECT  2.265 2.640 2.570 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.415 2.990 3.740 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.730 -0.180 1.540 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 0.840 1.525 1.180 ;
        RECT  1.185 0.840 1.525 1.685 ;
        RECT  1.185 1.455 2.035 1.685 ;
        RECT  1.770 1.455 2.035 3.170 ;
        RECT  0.810 2.940 2.035 3.170 ;
        RECT  0.810 2.940 1.150 3.450 ;
        RECT  1.960 0.565 3.740 0.870 ;
        RECT  1.960 0.470 2.300 1.225 ;
    END
END NAND2_A_OAI21_X2_18_SVT_WB

MACRO NAND2_A_OAI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_OAI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.415 2.330 0.980 2.730 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.685 1.540 2.260 ;
        RECT  1.010 1.685 1.540 1.965 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.365 1.720 2.705 2.260 ;
        RECT  2.255 1.720 2.705 2.040 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.470 1.770 3.780 2.425 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.385 2.960 3.220 3.300 ;
        RECT  2.935 1.015 3.220 3.300 ;
        RECT  2.760 1.015 3.220 1.355 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.170 2.960 0.535 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.400 -0.180 1.740 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.175 0.860 0.610 1.200 ;
        RECT  0.175 0.915 2.025 1.200 ;
        RECT  1.795 0.915 2.025 3.300 ;
        RECT  1.795 2.390 2.155 3.300 ;
        RECT  0.940 2.960 2.155 3.300 ;
    END
END NAND2_A_OAI21_X1_18_SVT_WB

MACRO NAND2_A_OAI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_OAI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.220 0.745 2.775 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.770 1.540 2.450 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.365 1.730 2.705 2.330 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.395 2.140 3.780 2.810 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.935 1.100 3.250 1.635 ;
        RECT  2.365 2.820 3.165 3.050 ;
        RECT  2.935 1.100 3.165 3.050 ;
        RECT  2.760 1.100 3.250 1.440 ;
        RECT  2.365 2.820 2.670 3.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.170 3.045 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.860 -0.180 1.670 0.480 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 0.980 2.135 1.320 ;
        RECT  1.845 0.980 2.135 3.050 ;
        RECT  0.975 2.820 2.135 3.050 ;
        RECT  0.975 2.820 1.280 3.330 ;
    END
END NAND2_A_OAI21_X0_18_SVT_WB

MACRO NAND2_A_NOR3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NOR3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.620 1.540 2.150 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.620 0.750 2.210 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.580 1.455 4.920 1.905 ;
        RECT  2.785 1.455 4.920 1.685 ;
        RECT  2.785 1.455 3.270 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.560 2.135 4.900 2.710 ;
        RECT  3.860 2.135 4.900 2.365 ;
        RECT  3.860 1.915 4.200 2.365 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.479  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 0.995 5.460 1.225 ;
        RECT  5.080 0.470 5.460 1.225 ;
        RECT  3.300 2.595 3.980 2.825 ;
        RECT  3.640 0.485 3.980 1.225 ;
        RECT  3.300 2.330 3.630 2.825 ;
        RECT  2.325 2.330 3.630 2.575 ;
        RECT  2.325 0.995 2.555 2.575 ;
        RECT  2.230 0.525 2.540 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.610 2.410 5.895 4.100 ;
        RECT  1.660 3.515 2.000 4.100 ;
        RECT  0.180 2.640 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.360 -0.180 4.700 0.765 ;
        RECT  2.920 -0.180 3.260 0.765 ;
        RECT  1.330 -0.180 1.670 0.930 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.650 0.520 1.390 ;
        RECT  0.180 1.160 2.000 1.390 ;
        RECT  1.770 1.160 2.000 3.285 ;
        RECT  5.150 1.840 5.640 2.180 ;
        RECT  1.770 1.840 2.095 3.285 ;
        RECT  0.900 2.575 2.095 3.285 ;
        RECT  5.150 1.840 5.380 3.285 ;
        RECT  0.900 3.055 5.380 3.285 ;
        RECT  0.900 2.575 1.240 3.385 ;
    END
END NAND2_A_NOR3_X4_18_SVT_WB

MACRO NAND2_A_NOR3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NOR3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.985 2.375 1.565 2.710 ;
        RECT  1.260 1.900 1.565 2.710 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.670 0.755 2.375 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.620 3.260 2.570 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.490 1.620 3.875 2.165 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.623  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.830 2.435 4.340 3.135 ;
        RECT  4.105 0.650 4.340 3.135 ;
        RECT  2.440 1.160 4.340 1.390 ;
        RECT  3.960 0.650 4.340 1.390 ;
        RECT  2.440 0.685 2.780 1.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  2.025 3.430 2.310 4.100 ;
        RECT  0.330 2.955 0.670 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.200 -0.180 3.540 0.930 ;
        RECT  1.680 -0.180 2.020 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.370 1.100 0.710 1.440 ;
        RECT  0.370 1.200 2.135 1.440 ;
        RECT  1.795 1.200 2.135 2.180 ;
        RECT  1.795 1.840 2.540 2.180 ;
        RECT  1.795 1.200 2.025 3.170 ;
        RECT  1.090 2.940 2.025 3.170 ;
        RECT  1.090 2.940 1.430 3.450 ;
    END
END NAND2_A_NOR3_X2_18_SVT_WB

MACRO NAND2_A_NOR3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NOR3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 2.070 1.580 2.865 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.025 0.900 2.305 ;
        RECT  0.140 2.025 0.690 2.835 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.325 1.600 2.710 2.100 ;
        RECT  2.325 1.430 2.630 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.535 3.325 2.345 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.811  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.480 2.620 3.785 3.270 ;
        RECT  3.555 0.860 3.785 3.270 ;
        RECT  2.050 0.860 3.785 1.200 ;
        RECT  3.200 2.620 3.785 2.960 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.180 3.095 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.635 -0.180 2.805 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.910 0.520 1.795 ;
        RECT  0.180 1.565 2.095 1.795 ;
        RECT  1.810 1.565 2.095 3.325 ;
        RECT  0.900 3.095 2.095 3.325 ;
        RECT  0.900 3.095 1.240 3.435 ;
    END
END NAND2_A_NOR3_X1_18_SVT_WB

MACRO NAND2_A_NOR3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NOR3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.880 1.440 2.170 ;
        RECT  0.140 1.880 0.570 2.710 ;
        END
    END AN
    PIN BN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.270 1.190 1.005 1.600 ;
        END
    END BN
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.375 1.410 2.830 1.750 ;
        RECT  2.375 1.410 2.660 2.150 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 2.080 3.270 2.870 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.400 3.070 3.780 3.410 ;
        RECT  3.500 0.890 3.780 3.410 ;
        RECT  3.170 0.890 3.780 1.250 ;
        RECT  2.010 0.890 3.780 1.180 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.180 3.515 1.880 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.595 -0.180 2.765 0.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.470 0.530 0.950 ;
        RECT  0.190 0.720 1.780 0.950 ;
        RECT  1.550 0.720 1.780 1.660 ;
        RECT  1.550 1.410 2.055 1.660 ;
        RECT  1.795 1.410 2.055 2.740 ;
        RECT  0.860 2.400 2.055 2.740 ;
    END
END NAND2_A_NOR3_X0_18_SVT_WB

MACRO NAND2_A_NAND2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NAND2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.640 1.745 1.040 2.250 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.420 1.260 1.760 1.980 ;
        RECT  1.210 1.260 1.760 1.585 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.635 3.750 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.809  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.460 2.940 4.925 3.170 ;
        RECT  4.610 1.160 4.925 3.170 ;
        RECT  3.180 1.160 4.925 1.405 ;
        RECT  3.850 2.940 4.190 3.450 ;
        RECT  3.180 0.685 3.520 1.405 ;
        RECT  2.460 2.940 2.800 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  1.700 3.045 2.040 4.100 ;
        RECT  0.170 2.545 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.370 -0.180 4.710 0.930 ;
        RECT  1.700 -0.180 2.040 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 0.580 2.580 0.880 ;
        RECT  0.220 0.580 0.560 1.360 ;
        RECT  2.240 0.580 2.580 2.710 ;
        RECT  2.240 2.380 4.380 2.710 ;
        RECT  4.090 1.860 4.380 2.710 ;
        RECT  0.940 2.480 4.380 2.710 ;
        RECT  0.940 2.480 1.280 3.235 ;
    END
END NAND2_A_NAND2_X4_18_SVT_WB

MACRO NAND2_A_NAND2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NAND2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.660 0.800 2.220 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 2.215 1.540 2.710 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.810 1.770 3.220 2.370 ;
        RECT  2.810 1.620 3.095 2.370 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.167  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.275 1.090 3.220 1.390 ;
        RECT  2.690 0.630 3.220 1.390 ;
        RECT  2.275 2.600 2.680 3.445 ;
        RECT  2.275 1.090 2.580 3.445 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 2.955 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.540 -0.180 1.880 0.905 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.090 0.560 1.430 ;
        RECT  0.220 1.200 2.045 1.430 ;
        RECT  1.790 1.200 2.045 3.170 ;
        RECT  0.940 2.940 2.045 3.170 ;
        RECT  0.940 2.940 1.280 3.450 ;
    END
END NAND2_A_NAND2_X2_18_SVT_WB

MACRO NAND2_A_NAND2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NAND2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.710 0.915 2.185 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.155 1.965 1.540 2.725 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.820 2.740 2.575 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.562  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.940 3.220 3.295 ;
        RECT  2.970 0.855 3.220 3.295 ;
        RECT  2.820 2.805 3.220 3.295 ;
        RECT  2.695 0.855 3.220 1.195 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.220 3.010 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.505 -0.180 1.845 0.820 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.855 0.520 1.340 ;
        RECT  0.180 1.110 2.070 1.340 ;
        RECT  1.785 1.110 2.070 3.295 ;
        RECT  0.940 2.955 2.070 3.295 ;
    END
END NAND2_A_NAND2_X1_18_SVT_WB

MACRO NAND2_A_NAND2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2_A_NAND2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.820 1.030 2.100 ;
        RECT  0.420 1.820 0.760 2.380 ;
        END
    END A0N
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.145 2.315 1.540 2.850 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 1.770 2.680 2.220 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 3.080 3.245 3.420 ;
        RECT  2.910 1.160 3.245 3.420 ;
        RECT  2.480 1.160 3.245 1.500 ;
        RECT  2.480 0.715 2.820 1.500 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 3.080 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.330 -0.180 1.670 1.055 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.715 0.520 1.590 ;
        RECT  0.180 1.285 2.000 1.590 ;
        RECT  1.770 2.510 2.150 2.850 ;
        RECT  1.770 1.285 2.000 3.420 ;
        RECT  0.900 3.080 2.000 3.420 ;
    END
END NAND2_A_NAND2_X0_18_SVT_WB

MACRO NAND2T_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.800 1.620 5.855 2.160 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.205 1.640 7.525 2.185 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.618  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.190 2.420 8.735 3.175 ;
        RECT  6.750 1.075 8.550 1.410 ;
        RECT  7.905 1.075 8.270 2.660 ;
        RECT  3.915 2.420 8.735 2.660 ;
        RECT  6.750 2.420 7.090 3.175 ;
        RECT  5.275 2.420 5.650 3.220 ;
        RECT  3.915 2.420 4.210 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  8.965 2.640 9.195 4.100 ;
        RECT  7.470 2.945 7.810 4.100 ;
        RECT  6.030 3.110 6.370 4.100 ;
        RECT  4.590 2.890 4.900 4.100 ;
        RECT  3.150 2.420 3.490 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  5.310 -0.180 5.650 0.800 ;
        RECT  3.870 -0.180 4.210 0.900 ;
        RECT  2.430 -0.180 2.770 0.900 ;
        RECT  0.990 -0.180 1.330 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  6.030 0.560 9.250 0.845 ;
        RECT  4.590 0.615 4.930 1.370 ;
        RECT  0.270 0.615 0.610 1.370 ;
        RECT  1.710 0.615 2.050 1.370 ;
        RECT  3.150 0.615 3.490 1.370 ;
        RECT  4.590 1.120 6.370 1.370 ;
        RECT  6.030 0.560 6.370 1.370 ;
        RECT  0.270 1.130 6.370 1.370 ;
        RECT  8.965 0.560 9.250 1.375 ;
    END
END NAND2T_X8_18_SVT_WB

MACRO NAND2T_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.245 1.600 5.030 2.210 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.715  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.830 1.680 3.635 2.300 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.126  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.745 1.105 6.525 1.345 ;
        RECT  6.185 0.590 6.525 1.345 ;
        RECT  5.465 2.530 6.020 3.395 ;
        RECT  5.700 1.105 6.020 3.395 ;
        RECT  4.000 2.530 6.020 2.810 ;
        RECT  4.745 1.005 5.085 1.345 ;
        RECT  4.000 2.530 4.365 3.340 ;
        RECT  0.905 2.530 6.020 2.760 ;
        RECT  2.400 2.530 2.690 3.340 ;
        RECT  0.905 2.530 1.245 3.315 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  6.250 2.630 6.535 4.100 ;
        RECT  4.745 3.165 5.085 4.100 ;
        RECT  3.065 3.075 3.405 4.100 ;
        RECT  1.625 3.090 1.965 4.100 ;
        RECT  0.180 2.990 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  3.065 -0.180 3.405 0.820 ;
        RECT  1.620 -0.180 1.960 0.820 ;
        RECT  0.180 -0.180 0.520 0.820 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  4.025 0.535 5.805 0.775 ;
        RECT  5.465 0.535 5.805 0.875 ;
        RECT  0.895 0.590 1.240 1.345 ;
        RECT  2.340 0.590 2.680 1.345 ;
        RECT  0.895 1.050 2.680 1.345 ;
        RECT  4.025 0.535 4.365 1.345 ;
        RECT  0.895 1.070 4.365 1.345 ;
    END
END NAND2T_X6_18_SVT_WB

MACRO NAND2T_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.820 1.120 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.170  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.640 2.150 2.175 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.809  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 3.045 2.760 3.330 ;
        RECT  2.380 1.105 2.760 3.330 ;
        RECT  0.900 1.105 2.760 1.410 ;
        RECT  0.900 2.630 1.240 3.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  3.140 2.575 3.480 4.100 ;
        RECT  1.660 3.560 2.000 4.100 ;
        RECT  0.180 2.630 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  3.900 -0.180 4.240 0.405 ;
        RECT  2.380 -0.180 2.720 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.645 5.000 0.875 ;
        RECT  0.180 0.645 0.520 1.400 ;
        RECT  3.140 0.645 3.480 1.400 ;
        RECT  4.660 0.645 5.000 1.400 ;
    END
END NAND2T_X4_18_SVT_WB

MACRO NAND2T_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.830 1.455 2.150 2.205 ;
        RECT  1.685 1.455 2.150 2.140 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.585  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.560 1.455 1.455 2.205 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.125  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.535 2.435 2.705 2.665 ;
        RECT  2.380 0.470 2.705 2.665 ;
        RECT  1.535 2.435 1.875 3.360 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.255 3.075 2.595 4.100 ;
        RECT  0.815 2.440 1.155 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.925 -0.180 1.265 0.765 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.205 0.470 0.545 1.225 ;
        RECT  1.645 0.470 1.985 1.225 ;
        RECT  0.205 0.995 1.985 1.225 ;
    END
END NAND2T_X2_18_SVT_WB

MACRO NAND2T_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.310 1.590 2.430 ;
        RECT  1.115 1.310 1.590 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.292  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.555 1.820 1.030 2.430 ;
        RECT  0.555 1.600 0.885 2.430 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.562  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.995 2.660 2.100 2.890 ;
        RECT  1.820 0.575 2.100 2.890 ;
        RECT  1.635 0.575 2.100 0.915 ;
        RECT  0.995 2.660 1.335 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.720 3.120 2.060 4.100 ;
        RECT  0.235 2.990 0.575 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.315 -0.180 0.655 1.330 ;
        END
    END VSS
END NAND2T_X1_18_SVT_WB

MACRO NAND2T_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.168  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.475 1.640 14.110 2.185 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.662  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.775 9.125 2.460 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.356  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.580 1.160 15.160 2.855 ;
        RECT  14.340 2.420 14.680 3.230 ;
        RECT  10.020 1.075 14.680 1.410 ;
        RECT  10.020 2.420 15.160 2.660 ;
        RECT  12.900 2.420 13.240 3.230 ;
        RECT  11.440 2.420 11.815 3.225 ;
        RECT  10.020 2.420 10.360 3.175 ;
        RECT  0.180 2.690 10.360 2.920 ;
        RECT  8.580 2.690 8.920 3.230 ;
        RECT  7.140 2.690 7.480 3.230 ;
        RECT  5.700 2.690 6.040 3.235 ;
        RECT  4.260 2.690 4.600 3.235 ;
        RECT  2.820 2.690 3.160 3.230 ;
        RECT  1.500 2.690 1.840 3.230 ;
        RECT  0.180 2.690 0.520 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  15.060 3.110 15.400 4.100 ;
        RECT  13.620 3.130 13.960 4.100 ;
        RECT  12.235 3.110 12.465 4.100 ;
        RECT  10.740 2.945 11.080 4.100 ;
        RECT  9.300 3.160 9.640 4.100 ;
        RECT  7.860 3.155 8.205 4.100 ;
        RECT  6.420 3.160 6.760 4.100 ;
        RECT  4.980 3.160 5.320 4.100 ;
        RECT  3.540 3.160 3.880 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  8.580 -0.180 8.920 0.800 ;
        RECT  7.140 -0.180 7.480 0.900 ;
        RECT  4.380 -0.180 4.720 0.900 ;
        RECT  2.940 -0.180 3.280 0.840 ;
        RECT  0.180 -0.180 0.520 0.845 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  9.300 0.555 15.400 0.845 ;
        RECT  15.060 0.555 15.400 0.905 ;
        RECT  7.860 0.615 8.200 1.365 ;
        RECT  3.660 0.615 4.000 1.365 ;
        RECT  5.100 0.615 5.440 1.365 ;
        RECT  6.420 0.615 6.760 1.365 ;
        RECT  0.900 0.560 1.240 1.365 ;
        RECT  2.220 0.560 2.560 1.365 ;
        RECT  7.860 1.120 9.640 1.365 ;
        RECT  3.660 1.130 9.640 1.365 ;
        RECT  9.300 0.555 9.640 1.365 ;
        RECT  0.900 1.135 9.640 1.365 ;
    END
END NAND2T_X16_18_SVT_WB

MACRO NAND2T_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.555 1.640 10.745 2.185 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.315  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.735 1.775 7.205 2.460 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.220 1.255 11.775 2.845 ;
        RECT  8.100 1.075 11.465 1.410 ;
        RECT  10.980 2.420 11.320 3.230 ;
        RECT  8.100 2.420 11.775 2.660 ;
        RECT  9.520 2.420 9.895 3.225 ;
        RECT  8.100 2.420 8.440 3.175 ;
        RECT  0.900 2.690 8.440 2.920 ;
        RECT  6.660 2.690 7.000 3.230 ;
        RECT  5.220 2.690 5.560 3.230 ;
        RECT  3.780 2.690 4.120 3.235 ;
        RECT  2.340 2.690 2.680 3.235 ;
        RECT  0.900 2.690 1.240 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.720 3.105 12.060 4.100 ;
        RECT  10.315 3.110 10.545 4.100 ;
        RECT  8.820 2.945 9.160 4.100 ;
        RECT  7.380 3.160 7.720 4.100 ;
        RECT  5.940 3.155 6.285 4.100 ;
        RECT  4.500 3.160 4.840 4.100 ;
        RECT  3.060 3.160 3.400 4.100 ;
        RECT  1.620 3.160 1.960 4.100 ;
        RECT  0.180 3.115 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  6.660 -0.180 7.000 0.800 ;
        RECT  5.220 -0.180 5.560 0.900 ;
        RECT  3.780 -0.180 4.120 0.900 ;
        RECT  2.340 -0.180 2.680 0.900 ;
        RECT  0.900 -0.180 1.240 0.840 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  7.380 0.555 12.040 0.845 ;
        RECT  11.700 0.555 12.040 0.940 ;
        RECT  5.940 0.615 6.280 1.365 ;
        RECT  1.620 0.615 1.960 1.365 ;
        RECT  3.060 0.615 3.400 1.365 ;
        RECT  4.500 0.615 4.840 1.365 ;
        RECT  0.180 0.560 0.520 1.365 ;
        RECT  5.940 1.120 7.720 1.365 ;
        RECT  1.620 1.130 7.720 1.365 ;
        RECT  7.380 0.555 7.720 1.365 ;
        RECT  0.180 1.135 7.720 1.365 ;
    END
END NAND2T_X12_18_SVT_WB

MACRO NAND2T_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN NAND2T_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.230 1.825 1.590 2.340 ;
        RECT  1.260 1.530 1.590 2.340 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.260 1.030 1.590 ;
        RECT  0.540 1.260 0.875 2.340 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.040 2.670 2.100 3.220 ;
        RECT  1.820 1.010 2.100 3.220 ;
        RECT  1.605 1.010 2.100 1.295 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.280 3.505 2.050 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.280 -0.180 0.620 1.030 ;
        END
    END VSS
END NAND2T_X0_18_SVT_WB

MACRO MUXI2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.695 4.470 2.190 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.235 1.770 1.580 2.360 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.770 2.380 8.110 3.190 ;
        RECT  6.450 1.050 8.110 1.390 ;
        RECT  7.770 0.580 8.110 1.390 ;
        RECT  7.420 1.050 7.770 2.655 ;
        RECT  6.450 2.380 8.110 2.655 ;
        RECT  6.450 2.380 6.790 3.190 ;
        RECT  6.450 0.580 6.790 1.390 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.260 2.865 1.980 ;
        RECT  0.575 1.260 2.865 1.540 ;
        RECT  0.575 1.260 0.860 1.655 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  4.410 2.420 4.750 4.100 ;
        RECT  0.960 3.515 1.300 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  4.410 -0.180 4.750 0.810 ;
        RECT  1.000 -0.180 1.340 1.030 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.690 0.620 1.030 ;
        RECT  0.115 0.690 0.345 3.180 ;
        RECT  1.910 1.860 2.215 3.180 ;
        RECT  0.115 2.830 2.215 3.180 ;
        RECT  3.555 1.630 3.830 3.180 ;
        RECT  0.115 2.950 3.830 3.180 ;
        RECT  3.095 1.060 4.930 1.400 ;
        RECT  4.700 1.060 4.930 2.185 ;
        RECT  4.700 1.845 5.690 2.185 ;
        RECT  3.095 1.060 3.325 2.720 ;
        RECT  2.445 2.380 3.325 2.720 ;
        RECT  5.160 0.470 5.470 1.280 ;
        RECT  5.160 0.940 6.220 1.280 ;
        RECT  5.990 1.620 6.550 1.960 ;
        RECT  5.990 0.940 6.220 2.760 ;
        RECT  5.130 2.420 6.220 2.760 ;
        RECT  5.130 2.420 5.470 3.230 ;
    END
END MUXI2_X8_18_SVT_WB

MACRO MUXI2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.355 1.770 3.830 2.380 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.135 1.100 1.595 1.540 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.320 2.235 7.660 3.410 ;
        RECT  6.000 1.145 7.660 1.440 ;
        RECT  7.320 0.535 7.660 1.440 ;
        RECT  6.000 2.235 7.660 2.465 ;
        RECT  6.795 1.145 7.260 2.465 ;
        RECT  6.000 2.235 6.340 3.385 ;
        RECT  6.000 0.535 6.340 1.440 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.695 1.770 2.205 2.000 ;
        RECT  1.920 1.570 2.205 2.000 ;
        RECT  0.695 1.770 1.035 2.150 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.240 3.030 5.580 4.100 ;
        RECT  3.780 2.880 4.120 4.100 ;
        RECT  0.970 3.515 1.310 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.240 -0.180 5.580 0.970 ;
        RECT  3.815 -0.180 4.120 0.915 ;
        RECT  0.930 -0.180 1.270 0.870 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.210 0.575 0.550 0.915 ;
        RECT  1.700 2.240 2.205 2.580 ;
        RECT  0.210 0.575 0.465 3.100 ;
        RECT  0.210 2.760 1.930 3.100 ;
        RECT  1.700 2.240 1.930 3.510 ;
        RECT  1.590 2.760 1.930 3.510 ;
        RECT  2.895 1.095 3.125 3.510 ;
        RECT  1.590 3.280 3.125 3.510 ;
        RECT  2.360 0.525 3.585 0.865 ;
        RECT  3.355 0.525 3.585 1.430 ;
        RECT  3.355 1.200 4.305 1.430 ;
        RECT  4.060 1.200 4.305 2.180 ;
        RECT  4.060 1.840 5.045 2.180 ;
        RECT  2.435 0.525 2.665 3.050 ;
        RECT  2.160 2.810 2.665 3.050 ;
        RECT  4.535 0.535 4.820 1.610 ;
        RECT  4.535 1.380 5.770 1.610 ;
        RECT  5.430 1.380 5.770 2.750 ;
        RECT  4.480 2.410 5.770 2.750 ;
        RECT  4.480 2.410 4.820 3.385 ;
    END
END MUXI2_X6_18_SVT_WB

MACRO MUXI2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 2.040 3.805 2.710 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.100 1.670 1.540 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.165 0.535 6.580 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.770 2.350 2.000 ;
        RECT  2.010 1.450 2.350 2.000 ;
        RECT  0.700 1.770 1.200 2.150 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.405 3.010 5.745 4.100 ;
        RECT  3.945 2.900 4.285 4.100 ;
        RECT  1.060 3.515 1.400 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  5.405 -0.180 5.745 0.970 ;
        RECT  3.960 -0.180 4.285 0.920 ;
        RECT  1.100 -0.180 1.440 0.870 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.240 0.580 0.720 0.920 ;
        RECT  1.790 2.230 2.350 2.525 ;
        RECT  0.240 0.580 0.470 3.060 ;
        RECT  0.240 2.720 2.020 3.060 ;
        RECT  1.790 2.230 2.020 3.510 ;
        RECT  1.680 2.720 2.020 3.510 ;
        RECT  3.040 1.100 3.270 3.510 ;
        RECT  1.680 3.280 3.270 3.510 ;
        RECT  2.480 0.530 3.730 0.870 ;
        RECT  3.500 0.530 3.730 1.810 ;
        RECT  3.500 1.470 4.415 1.810 ;
        RECT  4.160 1.470 4.415 2.175 ;
        RECT  4.160 1.820 5.260 2.175 ;
        RECT  2.580 0.530 2.810 3.050 ;
        RECT  2.250 2.755 2.810 3.050 ;
        RECT  4.645 0.535 4.985 1.440 ;
        RECT  4.645 1.210 5.935 1.440 ;
        RECT  5.595 1.210 5.935 2.745 ;
        RECT  4.645 2.405 5.935 2.745 ;
        RECT  4.645 2.405 4.985 3.385 ;
    END
END MUXI2_X4_18_SVT_WB

MACRO MUXI2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.770 3.840 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.100 1.670 1.540 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.891  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.145 0.535 6.580 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.770 2.350 2.000 ;
        RECT  2.010 1.445 2.350 2.000 ;
        RECT  0.700 1.770 1.200 2.155 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.385 3.050 5.725 4.100 ;
        RECT  3.925 2.870 4.265 4.100 ;
        RECT  1.060 3.515 1.400 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  5.385 -0.180 5.725 0.970 ;
        RECT  3.960 -0.180 4.265 0.925 ;
        RECT  1.100 -0.180 1.440 0.870 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.240 0.585 0.720 0.925 ;
        RECT  1.790 2.230 2.350 2.525 ;
        RECT  0.240 0.585 0.470 3.055 ;
        RECT  0.240 2.715 2.020 3.055 ;
        RECT  1.790 2.230 2.020 3.510 ;
        RECT  1.680 2.715 2.020 3.510 ;
        RECT  3.040 1.105 3.270 3.510 ;
        RECT  1.680 3.280 3.270 3.510 ;
        RECT  2.480 0.535 3.730 0.875 ;
        RECT  3.500 0.535 3.730 1.540 ;
        RECT  3.500 1.200 4.395 1.540 ;
        RECT  4.070 1.200 4.395 2.180 ;
        RECT  4.070 1.840 5.260 2.180 ;
        RECT  2.580 0.535 2.810 3.050 ;
        RECT  2.250 2.755 2.810 3.050 ;
        RECT  4.625 0.535 4.965 1.610 ;
        RECT  4.625 1.380 5.915 1.610 ;
        RECT  5.575 1.380 5.915 2.750 ;
        RECT  4.625 2.410 5.915 2.750 ;
        RECT  4.625 2.410 4.965 3.385 ;
    END
END MUXI2_X3_18_SVT_WB

MACRO MUXI2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.640 4.530 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.830 1.590 2.660 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.913  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.425 2.380 3.345 2.720 ;
        RECT  3.105 0.630 3.345 2.720 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.260 2.875 1.960 ;
        RECT  0.575 1.260 2.875 1.600 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.430 2.440 4.770 4.100 ;
        RECT  0.960 3.515 1.300 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.430 -0.180 4.770 1.410 ;
        RECT  1.000 -0.180 1.340 0.975 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.690 0.620 1.030 ;
        RECT  0.115 0.690 0.345 3.230 ;
        RECT  1.910 1.860 2.195 3.230 ;
        RECT  0.115 2.890 2.195 3.230 ;
        RECT  3.575 1.860 3.830 3.230 ;
        RECT  0.115 3.000 3.830 3.230 ;
    END
END MUXI2_X2_18_SVT_WB

MACRO MUXI2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.420 1.595 3.785 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.755 1.745 2.175 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.030 2.940 3.190 3.280 ;
        RECT  2.960 0.470 3.190 3.280 ;
        RECT  2.210 0.470 3.190 0.810 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.975 1.295 2.255 2.090 ;
        RECT  0.800 1.295 2.255 1.525 ;
        RECT  0.575 1.760 1.030 2.100 ;
        RECT  0.800 1.295 1.030 2.100 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.220 3.510 3.560 4.100 ;
        RECT  0.840 3.515 1.180 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.420 -0.180 3.740 0.490 ;
        RECT  1.020 -0.180 1.360 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.995 0.570 1.335 ;
        RECT  0.115 0.995 0.345 2.710 ;
        RECT  2.485 1.095 2.730 2.710 ;
        RECT  0.115 2.420 2.730 2.710 ;
    END
END MUXI2_X1_18_SVT_WB

MACRO MUXI2_X1P5_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X1P5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.975 1.595 4.340 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.770 1.750 2.190 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.300 2.940 3.470 3.295 ;
        RECT  3.240 0.470 3.470 3.295 ;
        RECT  2.490 0.470 3.470 0.810 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.373  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 1.310 2.420 1.965 ;
        RECT  0.800 1.310 2.420 1.540 ;
        RECT  0.690 1.640 1.030 2.150 ;
        RECT  0.800 1.310 1.030 2.150 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.700 2.960 4.000 4.100 ;
        RECT  0.940 3.010 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.810 -0.180 4.150 1.330 ;
        RECT  1.130 -0.180 1.470 0.860 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 0.570 1.440 ;
        RECT  0.180 1.100 0.460 2.710 ;
        RECT  2.725 1.095 3.010 2.710 ;
        RECT  0.180 2.420 3.010 2.710 ;
    END
END MUXI2_X1P5_18_SVT_WB

MACRO MUXI2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.015 1.705 4.480 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.775 1.650 2.450 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.210 2.420 9.550 3.230 ;
        RECT  6.450 1.085 9.550 1.325 ;
        RECT  9.210 0.515 9.550 1.325 ;
        RECT  6.450 2.420 9.550 2.760 ;
        RECT  7.755 1.085 8.420 2.760 ;
        RECT  7.770 0.470 8.110 3.230 ;
        RECT  6.450 0.985 8.110 1.325 ;
        RECT  6.450 2.420 6.790 3.230 ;
        RECT  6.450 0.515 6.790 1.325 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.240 2.865 1.980 ;
        RECT  0.575 1.240 2.865 1.545 ;
        RECT  0.575 1.240 0.860 1.730 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.930 2.640 10.270 4.100 ;
        RECT  8.490 3.110 8.830 4.100 ;
        RECT  4.410 2.430 4.750 4.100 ;
        RECT  0.960 3.515 1.300 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.930 -0.180 10.270 1.325 ;
        RECT  8.490 -0.180 8.830 0.855 ;
        RECT  4.410 -0.180 4.750 0.810 ;
        RECT  1.000 -0.180 1.340 0.850 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.525 0.620 0.865 ;
        RECT  0.115 0.525 0.345 3.230 ;
        RECT  1.910 1.860 2.215 3.230 ;
        RECT  0.115 2.890 2.215 3.230 ;
        RECT  3.555 1.640 3.785 3.230 ;
        RECT  0.115 2.950 3.785 3.230 ;
        RECT  3.095 1.100 4.940 1.410 ;
        RECT  4.710 1.100 4.940 2.200 ;
        RECT  4.710 1.860 5.695 2.200 ;
        RECT  3.095 1.100 3.325 2.720 ;
        RECT  2.445 2.380 3.325 2.720 ;
        RECT  5.170 0.470 5.470 1.280 ;
        RECT  5.170 0.940 6.220 1.280 ;
        RECT  5.990 1.620 6.550 1.960 ;
        RECT  5.990 0.940 6.220 2.770 ;
        RECT  5.130 2.430 6.220 2.770 ;
        RECT  5.130 2.430 5.470 3.240 ;
    END
END MUXI2_X12_18_SVT_WB

MACRO MUXI2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.210 3.840 1.995 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.090 1.660 1.540 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.538  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.155 2.805 2.660 3.050 ;
        RECT  2.430 0.575 2.660 3.050 ;
        RECT  2.320 0.575 2.660 1.030 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.770 2.200 2.000 ;
        RECT  1.915 1.565 2.200 2.000 ;
        RECT  0.700 1.770 1.205 2.150 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.745 2.755 4.085 4.100 ;
        RECT  0.875 3.515 1.215 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.745 -0.180 4.085 0.915 ;
        RECT  1.005 -0.180 1.345 0.860 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.240 0.575 0.625 0.915 ;
        RECT  1.695 2.235 2.200 2.575 ;
        RECT  0.240 0.575 0.470 3.095 ;
        RECT  0.240 2.755 1.925 3.095 ;
        RECT  1.695 2.235 1.925 3.510 ;
        RECT  1.585 2.755 1.925 3.510 ;
        RECT  2.890 1.135 3.175 3.510 ;
        RECT  1.585 3.280 3.175 3.510 ;
    END
END MUXI2_X0_18_SVT_WB

MACRO MUXI2PG_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2PG_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.553  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.770 1.455 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.553  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.635 1.635 10.430 2.040 ;
        RECT  9.070 1.915 10.045 2.200 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.375  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 3.185 7.405 3.470 ;
        RECT  5.610 0.470 7.390 0.755 ;
        RECT  0.750 0.470 7.390 0.700 ;
        RECT  0.130 0.690 4.120 0.755 ;
        RECT  0.130 2.950 2.480 3.285 ;
        RECT  0.130 0.690 0.975 0.920 ;
        RECT  0.130 0.690 0.470 3.285 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.210 8.925 1.735 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.635 2.900 11.975 4.100 ;
        RECT  10.195 3.000 10.535 4.100 ;
        RECT  8.750 3.185 9.090 4.100 ;
        RECT  1.700 3.515 2.040 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.635 -0.180 11.975 0.795 ;
        RECT  10.195 -0.180 10.535 0.740 ;
        RECT  0.180 -0.180 0.520 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.460 0.985 4.785 1.270 ;
        RECT  4.480 0.930 4.785 1.270 ;
        RECT  0.940 1.150 2.970 1.440 ;
        RECT  2.460 0.985 2.970 2.720 ;
        RECT  0.940 2.380 2.970 2.720 ;
        RECT  2.740 0.985 2.970 2.955 ;
        RECT  2.740 2.725 6.800 2.955 ;
        RECT  5.475 1.450 8.310 1.790 ;
        RECT  8.080 0.870 8.310 2.495 ;
        RECT  7.985 1.450 8.310 2.495 ;
        RECT  7.985 2.155 8.325 2.495 ;
        RECT  7.620 0.410 9.530 0.640 ;
        RECT  9.300 0.410 9.530 1.270 ;
        RECT  7.620 0.410 7.850 1.220 ;
        RECT  5.015 0.985 7.850 1.220 ;
        RECT  9.300 0.970 11.255 1.270 ;
        RECT  5.015 0.985 5.245 2.495 ;
        RECT  4.880 2.210 5.245 2.495 ;
        RECT  10.915 0.970 11.255 2.770 ;
        RECT  9.530 2.430 11.255 2.770 ;
    END
END MUXI2PG_X8_18_SVT_WB

MACRO MUXI2PG_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2PG_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.775 1.770 1.540 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.035 1.810 10.095 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.343  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.995 0.470 6.775 0.755 ;
        RECT  2.270 3.185 6.730 3.470 ;
        RECT  6.435 3.110 6.730 3.470 ;
        RECT  0.750 0.470 6.775 0.700 ;
        RECT  0.140 0.690 3.505 0.755 ;
        RECT  0.140 2.950 2.480 3.285 ;
        RECT  0.140 0.690 0.975 0.920 ;
        RECT  0.140 0.690 0.480 3.285 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.157  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.420 1.910 7.700 2.710 ;
        RECT  7.280 1.910 7.700 2.200 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  10.680 3.460 11.020 4.100 ;
        RECT  1.700 3.515 2.040 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  10.640 -0.180 10.980 0.810 ;
        RECT  9.200 -0.180 9.540 0.890 ;
        RECT  0.180 -0.180 0.520 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.460 0.985 4.170 1.270 ;
        RECT  3.865 0.930 4.170 1.270 ;
        RECT  0.940 1.150 2.970 1.440 ;
        RECT  2.460 0.985 2.970 2.720 ;
        RECT  0.940 2.380 2.970 2.720 ;
        RECT  2.740 0.985 2.970 2.955 ;
        RECT  5.715 2.615 6.055 2.955 ;
        RECT  2.740 2.725 6.055 2.955 ;
        RECT  7.780 0.880 8.215 1.680 ;
        RECT  4.860 1.450 8.215 1.680 ;
        RECT  4.860 1.450 5.145 1.790 ;
        RECT  7.930 0.880 8.215 2.940 ;
        RECT  7.195 0.410 8.805 0.650 ;
        RECT  7.195 0.410 7.535 1.220 ;
        RECT  4.400 0.985 7.535 1.220 ;
        RECT  8.480 1.120 10.260 1.440 ;
        RECT  8.480 0.410 8.805 2.720 ;
        RECT  4.400 0.985 4.630 2.495 ;
        RECT  4.265 2.210 4.630 2.495 ;
        RECT  8.480 2.380 10.260 2.720 ;
    END
END MUXI2PG_X6_18_SVT_WB

MACRO MUXI2PG_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2PG_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.670 0.990 2.250 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.765  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.325 2.100 2.470 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.350 2.230 6.285 2.515 ;
        RECT  6.055 0.700 6.285 2.515 ;
        RECT  5.350 0.700 6.285 1.290 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.575  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.470 3.675 1.760 ;
        RECT  2.940 1.080 3.280 1.760 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  1.665 3.560 2.005 4.100 ;
        RECT  0.185 2.630 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  1.665 -0.180 2.005 0.405 ;
        RECT  0.185 -0.180 0.525 1.290 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.865 1.005 4.245 1.290 ;
        RECT  3.970 1.520 5.825 1.860 ;
        RECT  3.970 1.005 4.245 2.515 ;
        RECT  3.905 2.230 4.245 2.515 ;
        RECT  2.425 0.470 4.970 0.775 ;
        RECT  2.425 0.470 2.700 2.815 ;
        RECT  2.425 2.475 2.935 2.815 ;
        RECT  2.705 2.745 6.410 2.975 ;
        RECT  0.905 0.590 1.245 1.345 ;
        RECT  6.515 0.480 6.800 2.515 ;
        RECT  1.220 1.115 1.450 3.330 ;
        RECT  0.905 2.630 1.450 3.330 ;
        RECT  0.905 3.045 2.485 3.330 ;
        RECT  6.745 2.175 7.085 3.510 ;
        RECT  2.235 3.205 7.085 3.510 ;
    END
END MUXI2PG_X4_18_SVT_WB

MACRO MUXI2D_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2D_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.265 3.805 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.640 2.780 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.563  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.915 2.410 9.320 3.380 ;
        RECT  7.595 1.265 9.320 1.550 ;
        RECT  8.915 0.530 9.320 1.550 ;
        RECT  7.595 2.405 8.945 2.660 ;
        RECT  8.365 1.265 8.945 2.660 ;
        RECT  7.595 2.405 7.975 3.385 ;
        RECT  7.595 0.535 7.975 1.550 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 2.705 5.405 2.935 ;
        RECT  5.170 1.860 5.405 2.935 ;
        RECT  1.140 2.950 5.115 3.285 ;
        RECT  4.520 2.705 5.115 3.285 ;
        RECT  1.140 1.640 1.480 3.285 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  6.835 3.515 7.175 4.100 ;
        RECT  5.355 3.165 5.695 4.100 ;
        RECT  1.370 3.515 1.710 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  6.835 -0.180 7.175 0.875 ;
        RECT  5.090 -0.180 5.430 0.890 ;
        RECT  0.900 -0.180 1.240 0.880 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.810 0.530 4.420 0.870 ;
        RECT  0.180 1.110 2.150 1.410 ;
        RECT  4.135 0.530 4.420 1.980 ;
        RECT  1.810 0.530 2.150 2.200 ;
        RECT  0.180 0.540 0.520 3.095 ;
        RECT  4.650 1.305 5.865 1.535 ;
        RECT  5.635 1.305 5.865 2.180 ;
        RECT  5.635 1.835 6.660 2.180 ;
        RECT  4.650 1.305 4.880 2.440 ;
        RECT  4.040 2.210 4.880 2.440 ;
        RECT  3.010 1.100 3.270 2.710 ;
        RECT  2.720 2.380 3.270 2.710 ;
        RECT  4.040 2.210 4.270 2.710 ;
        RECT  2.720 2.480 4.270 2.710 ;
        RECT  6.095 0.535 6.415 1.540 ;
        RECT  6.095 1.310 7.365 1.540 ;
        RECT  7.085 1.310 7.365 2.915 ;
        RECT  6.075 2.575 7.365 2.915 ;
        RECT  6.075 2.575 6.415 3.385 ;
    END
END MUXI2D_X8_18_SVT_WB

MACRO MUXI2D_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2D_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.580 1.760 3.270 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.665 2.240 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 0.535 6.580 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.425 3.335 2.765 ;
        RECT  0.700 1.175 1.040 2.765 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.440 3.515 5.780 4.100 ;
        RECT  4.025 2.945 4.320 4.100 ;
        RECT  0.990 3.100 1.330 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  5.440 -0.180 5.780 0.875 ;
        RECT  4.025 -0.180 4.320 0.915 ;
        RECT  0.950 -0.180 1.290 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.575 0.530 0.940 ;
        RECT  0.190 0.635 1.610 0.940 ;
        RECT  1.270 0.635 1.610 1.435 ;
        RECT  1.270 1.095 3.335 1.435 ;
        RECT  1.270 0.635 1.570 2.195 ;
        RECT  0.190 0.575 0.470 3.440 ;
        RECT  0.190 3.100 0.610 3.440 ;
        RECT  2.140 0.470 3.795 0.810 ;
        RECT  3.565 1.840 5.260 2.180 ;
        RECT  3.565 0.470 3.795 3.405 ;
        RECT  2.140 3.065 3.795 3.405 ;
        RECT  4.680 0.535 5.020 1.385 ;
        RECT  4.680 1.105 5.970 1.385 ;
        RECT  5.685 1.105 5.970 2.815 ;
        RECT  4.680 2.475 5.970 2.815 ;
        RECT  4.680 2.475 5.020 3.385 ;
    END
END MUXI2D_X4_18_SVT_WB

MACRO MUXI2D_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2D_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.275 3.875 2.160 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.640 2.780 2.150 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.740 2.380 3.270 2.720 ;
        RECT  3.010 1.100 3.270 2.720 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.785 1.840 5.125 2.720 ;
        RECT  1.155 2.950 4.785 3.285 ;
        RECT  4.445 2.380 4.785 3.285 ;
        RECT  1.155 1.640 1.495 3.285 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  5.025 3.110 5.365 4.100 ;
        RECT  1.370 3.515 1.710 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  5.060 -0.180 5.400 1.345 ;
        RECT  0.915 -0.180 1.255 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.825 0.530 4.455 0.870 ;
        RECT  0.195 1.040 2.150 1.380 ;
        RECT  4.110 0.530 4.455 1.960 ;
        RECT  1.825 0.530 2.150 2.200 ;
        RECT  0.195 0.470 0.535 3.295 ;
    END
END MUXI2D_X2_18_SVT_WB

MACRO MUXI2D_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2D_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.570 1.770 3.270 2.115 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.675 2.230 2.175 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.130 3.005 3.785 3.345 ;
        RECT  3.555 0.535 3.785 3.345 ;
        RECT  2.130 0.535 3.785 0.875 ;
        RECT  2.130 0.535 2.710 0.980 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.545 3.325 2.775 ;
        RECT  3.040 2.435 3.325 2.775 ;
        RECT  0.700 1.185 1.040 2.775 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  4.015 3.110 4.300 4.100 ;
        RECT  0.980 3.110 1.320 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  4.015 -0.180 4.300 0.820 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.585 0.520 0.950 ;
        RECT  0.180 0.635 1.610 0.950 ;
        RECT  1.270 0.635 1.610 1.445 ;
        RECT  3.040 1.105 3.325 1.445 ;
        RECT  1.270 1.210 3.325 1.445 ;
        RECT  1.270 0.635 1.560 2.315 ;
        RECT  0.180 0.585 0.460 3.450 ;
        RECT  0.180 3.110 0.600 3.450 ;
    END
END MUXI2D_X1_18_SVT_WB

MACRO MUXI2D_X1P5_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2D_X1P5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 2.195 3.220 2.535 ;
        RECT  2.905 1.095 3.220 2.535 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 1.210 2.675 1.665 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.765 2.740 3.050 ;
        RECT  1.770 0.575 2.705 0.980 ;
        RECT  1.770 0.575 2.000 3.050 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.571  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.915 1.770 1.540 2.150 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.910 2.515 4.195 4.100 ;
        RECT  0.795 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.960 -0.180 4.300 1.305 ;
        RECT  1.080 -0.180 1.420 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.450 1.860 3.820 2.200 ;
        RECT  0.360 1.100 0.685 2.720 ;
        RECT  0.360 2.380 1.540 2.720 ;
        RECT  1.310 2.380 1.540 3.510 ;
        RECT  3.450 1.860 3.680 3.510 ;
        RECT  1.310 3.280 3.680 3.510 ;
    END
END MUXI2D_X1P5_18_SVT_WB

MACRO MUXI2D_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUXI2D_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.480 1.700 3.345 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.650 2.220 2.100 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.070 2.890 3.805 3.270 ;
        RECT  3.575 0.540 3.805 3.270 ;
        RECT  2.150 0.540 3.805 0.835 ;
        RECT  2.150 0.540 2.490 0.880 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.330 3.345 2.660 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.920 2.890 1.260 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.960 -0.180 1.300 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.540 0.540 1.530 ;
        RECT  3.060 1.065 3.345 1.420 ;
        RECT  0.190 1.190 3.345 1.420 ;
        RECT  0.190 1.190 1.500 1.530 ;
        RECT  1.160 1.190 1.500 1.830 ;
        RECT  0.190 0.540 0.420 3.230 ;
        RECT  0.190 2.890 0.540 3.230 ;
    END
END MUXI2D_X0_18_SVT_WB

MACRO MUX2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.975 1.700 4.340 2.255 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.770 1.735 2.200 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.570 2.575 6.910 3.400 ;
        RECT  5.175 1.055 6.910 1.345 ;
        RECT  6.570 0.535 6.910 1.345 ;
        RECT  5.175 2.575 6.910 2.865 ;
        RECT  5.740 1.055 6.120 2.865 ;
        RECT  5.175 2.575 5.470 3.385 ;
        RECT  5.175 0.535 5.470 1.345 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.650 1.200 2.935 2.200 ;
        RECT  0.695 1.200 2.935 1.540 ;
        RECT  0.695 1.200 0.980 2.150 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  7.290 2.590 7.630 4.100 ;
        RECT  5.850 3.095 6.190 4.100 ;
        RECT  4.370 2.955 4.710 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  7.290 -0.180 7.630 1.345 ;
        RECT  5.850 -0.180 6.190 0.825 ;
        RECT  4.370 -0.180 4.710 0.915 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.050 0.465 2.840 ;
        RECT  1.980 1.860 2.320 2.840 ;
        RECT  3.320 1.635 3.605 2.840 ;
        RECT  0.180 2.500 3.605 2.840 ;
        RECT  3.080 0.470 3.420 0.865 ;
        RECT  3.165 0.470 3.420 1.375 ;
        RECT  3.165 1.145 4.945 1.375 ;
        RECT  4.660 1.145 4.945 2.715 ;
        RECT  3.835 2.485 4.945 2.715 ;
        RECT  3.835 2.485 4.085 3.300 ;
        RECT  2.220 3.070 4.085 3.300 ;
        RECT  2.220 3.070 2.560 3.450 ;
    END
END MUX2_X8_18_SVT_WB

MACRO MUX2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.120 3.370 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.190 1.540 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.605 2.235 6.020 3.235 ;
        RECT  4.165 1.615 6.020 1.845 ;
        RECT  5.605 0.630 6.020 1.845 ;
        RECT  4.165 2.235 6.020 2.465 ;
        RECT  5.010 1.615 5.350 2.465 ;
        RECT  4.165 2.235 4.505 3.235 ;
        RECT  4.165 0.535 4.505 1.845 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.820 2.250 2.105 ;
        RECT  1.790 1.765 2.250 2.105 ;
        RECT  0.730 1.820 1.070 2.205 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.885 2.695 5.225 4.100 ;
        RECT  3.405 3.515 3.745 4.100 ;
        RECT  0.985 3.515 1.325 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.885 -0.180 5.225 1.385 ;
        RECT  3.405 -0.180 3.745 0.405 ;
        RECT  0.985 -0.180 1.325 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.225 0.575 0.565 0.915 ;
        RECT  0.225 0.635 2.000 0.915 ;
        RECT  1.770 0.635 2.000 1.435 ;
        RECT  1.770 1.095 2.710 1.435 ;
        RECT  2.480 1.095 2.710 2.775 ;
        RECT  0.225 2.435 2.710 2.775 ;
        RECT  0.225 2.435 0.565 3.295 ;
        RECT  2.230 0.525 2.515 0.865 ;
        RECT  2.230 0.635 3.935 0.865 ;
        RECT  3.600 0.635 3.935 3.285 ;
        RECT  2.175 3.005 3.935 3.285 ;
        RECT  2.175 3.005 2.515 3.345 ;
    END
END MUX2_X6_18_SVT_WB

MACRO MUX2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.095 3.370 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.210 1.540 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 0.535 4.505 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.730 1.915 2.250 2.150 ;
        RECT  1.820 1.765 2.250 2.150 ;
        RECT  0.730 1.915 1.070 2.255 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.885 2.575 5.225 4.100 ;
        RECT  3.405 3.515 3.745 4.100 ;
        RECT  0.985 3.515 1.325 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.885 -0.180 5.225 1.345 ;
        RECT  3.405 -0.180 3.745 0.405 ;
        RECT  0.985 -0.180 1.325 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.225 0.575 0.565 0.915 ;
        RECT  0.225 0.635 2.000 0.915 ;
        RECT  1.770 0.635 2.000 1.435 ;
        RECT  1.770 1.095 2.710 1.435 ;
        RECT  1.950 2.435 2.710 2.775 ;
        RECT  2.480 1.095 2.710 2.775 ;
        RECT  0.225 2.545 2.710 2.775 ;
        RECT  0.225 2.545 0.565 3.295 ;
        RECT  2.230 0.525 2.515 0.865 ;
        RECT  2.230 0.635 3.830 0.865 ;
        RECT  3.600 0.635 3.830 3.285 ;
        RECT  2.175 3.005 3.830 3.285 ;
        RECT  2.175 3.005 2.515 3.345 ;
    END
END MUX2_X4_18_SVT_WB

MACRO MUX2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.095 3.350 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.210 1.440 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.894  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 0.535 4.460 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.820 2.240 2.160 ;
        RECT  1.880 1.765 2.240 2.160 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.880 2.920 5.220 4.100 ;
        RECT  3.360 3.515 3.700 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.880 -0.180 5.220 0.970 ;
        RECT  3.360 -0.180 3.700 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.575 0.510 0.915 ;
        RECT  0.180 0.635 1.900 0.915 ;
        RECT  1.670 0.635 1.900 1.435 ;
        RECT  1.670 1.095 2.710 1.435 ;
        RECT  2.470 1.095 2.710 2.775 ;
        RECT  0.180 2.435 2.710 2.775 ;
        RECT  0.180 2.435 0.510 3.295 ;
        RECT  2.130 0.525 2.470 0.865 ;
        RECT  2.130 0.635 3.830 0.865 ;
        RECT  3.580 0.635 3.830 3.285 ;
        RECT  2.130 3.005 3.830 3.285 ;
        RECT  2.130 3.005 2.470 3.345 ;
    END
END MUX2_X3_18_SVT_WB

MACRO MUX2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.095 3.780 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.210 1.840 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 0.535 4.900 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.915 2.660 2.150 ;
        RECT  2.300 1.765 2.660 2.150 ;
        RECT  1.060 1.915 1.400 2.255 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.760 3.515 4.100 4.100 ;
        RECT  1.340 3.515 1.680 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.760 -0.180 4.100 0.405 ;
        RECT  1.340 -0.180 1.680 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.580 0.575 0.920 0.915 ;
        RECT  0.580 0.635 2.300 0.915 ;
        RECT  2.070 0.635 2.300 1.435 ;
        RECT  2.070 1.095 3.120 1.435 ;
        RECT  2.310 2.435 3.120 2.780 ;
        RECT  2.890 1.095 3.120 2.780 ;
        RECT  0.580 2.550 3.120 2.780 ;
        RECT  0.580 2.550 0.920 3.295 ;
        RECT  2.530 0.525 2.870 0.865 ;
        RECT  2.530 0.635 4.290 0.865 ;
        RECT  4.010 0.635 4.290 3.285 ;
        RECT  2.530 3.010 4.290 3.285 ;
        RECT  2.530 3.010 2.870 3.350 ;
    END
END MUX2_X2_18_SVT_WB

MACRO MUX2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.095 3.780 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.210 1.840 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 0.535 4.900 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.915 2.660 2.150 ;
        RECT  2.300 1.765 2.660 2.150 ;
        RECT  1.060 1.915 1.400 2.255 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.760 3.515 4.100 4.100 ;
        RECT  1.340 3.515 1.680 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.760 -0.180 4.100 0.405 ;
        RECT  1.340 -0.180 1.680 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.580 0.575 0.920 0.915 ;
        RECT  0.580 0.635 2.300 0.915 ;
        RECT  2.070 0.635 2.300 1.435 ;
        RECT  2.070 1.095 3.120 1.435 ;
        RECT  2.310 2.435 3.120 2.780 ;
        RECT  2.890 1.095 3.120 2.780 ;
        RECT  0.580 2.550 3.120 2.780 ;
        RECT  0.580 2.550 0.920 3.295 ;
        RECT  2.530 0.525 2.870 0.865 ;
        RECT  2.530 0.635 4.290 0.865 ;
        RECT  4.010 0.635 4.290 3.285 ;
        RECT  2.530 3.010 4.290 3.285 ;
        RECT  2.530 3.010 2.870 3.350 ;
    END
END MUX2_X1_18_SVT_WB

MACRO MUX2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.040 1.645 4.405 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.770 1.730 2.200 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.820 2.575 8.160 3.385 ;
        RECT  5.225 1.005 8.160 1.345 ;
        RECT  7.820 0.535 8.160 1.345 ;
        RECT  5.225 2.575 8.160 2.915 ;
        RECT  6.460 1.005 7.140 2.915 ;
        RECT  6.500 0.470 6.840 3.450 ;
        RECT  5.225 2.575 5.520 3.385 ;
        RECT  5.225 0.535 5.520 1.345 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.700 1.200 3.040 2.200 ;
        RECT  0.745 1.200 3.040 1.540 ;
        RECT  0.745 1.200 1.030 2.200 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  4.420 3.045 4.760 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  4.420 -0.180 4.760 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.220 1.100 0.515 2.770 ;
        RECT  2.030 1.860 2.370 2.770 ;
        RECT  3.370 1.640 3.710 2.770 ;
        RECT  0.220 2.430 3.710 2.770 ;
        RECT  3.130 0.470 3.500 0.810 ;
        RECT  3.270 0.470 3.500 1.410 ;
        RECT  3.270 1.105 4.995 1.410 ;
        RECT  4.710 1.105 4.995 2.785 ;
        RECT  3.940 2.445 4.995 2.785 ;
        RECT  3.940 2.445 4.190 3.450 ;
        RECT  2.420 3.110 4.190 3.450 ;
    END
END MUX2_X12_18_SVT_WB

MACRO MUX2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN MUX2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.370 1.095 3.780 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.210 1.840 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 0.535 4.900 3.295 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.915 2.660 2.150 ;
        RECT  2.300 1.765 2.660 2.150 ;
        RECT  1.060 1.915 1.400 2.255 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.760 3.515 4.100 4.100 ;
        RECT  1.340 3.515 1.680 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.760 -0.180 4.100 0.405 ;
        RECT  1.340 -0.180 1.680 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.580 0.575 0.920 0.915 ;
        RECT  0.580 0.635 2.300 0.915 ;
        RECT  2.070 0.635 2.300 1.435 ;
        RECT  2.070 1.095 3.120 1.435 ;
        RECT  2.310 2.435 3.120 2.780 ;
        RECT  2.890 1.095 3.120 2.780 ;
        RECT  0.580 2.550 3.120 2.780 ;
        RECT  0.580 2.550 0.920 3.295 ;
        RECT  2.530 0.525 2.870 0.865 ;
        RECT  2.530 0.635 4.290 0.865 ;
        RECT  4.010 0.635 4.290 3.285 ;
        RECT  2.530 3.010 4.290 3.285 ;
        RECT  2.530 3.010 2.870 3.350 ;
    END
END MUX2_X0_18_SVT_WB

MACRO INV_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.615 1.665 1.565 2.160 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.570 2.560 3.390 ;
        RECT  0.900 0.955 2.560 1.295 ;
        RECT  2.220 0.470 2.560 1.295 ;
        RECT  0.900 2.570 2.560 2.920 ;
        RECT  1.795 0.955 2.160 2.920 ;
        RECT  0.900 2.570 1.240 3.390 ;
        RECT  0.900 0.475 1.240 1.295 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 2.580 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.180 -0.180 0.520 1.320 ;
        END
    END VSS
END INV_X8_18_SVT_WB

MACRO INV_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.620 1.565 2.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.380 2.560 3.190 ;
        RECT  0.900 1.015 2.560 1.290 ;
        RECT  2.220 0.480 2.560 1.290 ;
        RECT  0.900 2.380 2.560 2.660 ;
        RECT  1.795 1.015 2.105 2.660 ;
        RECT  0.900 2.380 1.240 3.190 ;
        RECT  0.900 0.480 1.240 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.600 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.180 -0.180 0.520 1.290 ;
        END
    END VSS
END INV_X6_18_SVT_WB

MACRO INV_X5_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.988  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.610 1.010 2.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.867  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.380 2.560 3.255 ;
        RECT  0.895 0.865 2.560 1.200 ;
        RECT  0.915 2.380 2.560 2.685 ;
        RECT  1.775 0.865 2.150 2.685 ;
        RECT  0.915 2.380 1.240 3.255 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.445 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.180 -0.180 0.520 0.985 ;
        END
    END VSS
END INV_X5_18_SVT_WB

MACRO INV_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.615 1.005 1.960 ;
        RECT  0.140 1.615 0.485 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.298  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.235 0.985 1.545 2.440 ;
        RECT  1.000 2.220 1.340 3.190 ;
        RECT  0.980 0.495 1.295 1.250 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.720 2.620 2.060 4.100 ;
        RECT  0.230 2.600 0.570 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.775 -0.180 2.060 1.320 ;
        RECT  0.230 -0.180 0.570 1.230 ;
        END
    END VSS
END INV_X4_18_SVT_WB

MACRO INV_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.260 1.590 1.795 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.888  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.905 2.405 1.245 2.915 ;
        RECT  0.700 0.650 1.245 1.030 ;
        RECT  0.700 0.650 0.930 2.635 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.625 2.820 1.965 4.100 ;
        RECT  0.185 2.820 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.625 -0.180 1.965 0.865 ;
        RECT  0.185 -0.180 0.470 0.865 ;
        END
    END VSS
END INV_X3_18_SVT_WB

MACRO INV_X32_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X32_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.940  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 1.620 6.450 2.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.372  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.240 2.400 11.580 3.390 ;
        RECT  1.145 0.990 11.580 1.255 ;
        RECT  11.240 0.470 11.580 1.255 ;
        RECT  1.210 2.400 11.580 2.740 ;
        RECT  9.800 2.400 10.140 3.390 ;
        RECT  9.800 0.470 10.140 1.255 ;
        RECT  8.360 2.400 8.700 3.210 ;
        RECT  8.360 0.470 8.700 1.255 ;
        RECT  6.920 2.400 8.700 2.745 ;
        RECT  6.850 0.990 7.595 2.740 ;
        RECT  6.920 0.470 7.260 3.230 ;
        RECT  5.480 2.400 5.820 3.230 ;
        RECT  5.480 0.470 5.820 1.255 ;
        RECT  4.040 2.400 4.380 3.230 ;
        RECT  4.040 0.470 4.380 1.255 ;
        RECT  2.600 2.400 2.940 3.230 ;
        RECT  2.600 0.470 2.940 1.255 ;
        RECT  1.210 2.400 2.940 2.745 ;
        RECT  1.210 2.400 1.500 3.230 ;
        RECT  1.145 0.470 1.500 1.255 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  10.520 3.100 10.860 4.100 ;
        RECT  9.080 3.100 9.420 4.100 ;
        RECT  7.640 3.155 7.980 4.100 ;
        RECT  6.200 3.160 6.540 4.100 ;
        RECT  4.760 3.155 5.100 4.100 ;
        RECT  3.320 3.150 3.660 4.100 ;
        RECT  1.880 3.140 2.220 4.100 ;
        RECT  0.440 2.640 0.780 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  10.520 -0.180 10.860 0.760 ;
        RECT  9.080 -0.180 9.420 0.760 ;
        RECT  7.640 -0.180 7.980 0.760 ;
        RECT  6.200 -0.180 6.540 0.760 ;
        RECT  4.760 -0.180 5.100 0.760 ;
        RECT  3.320 -0.180 3.660 0.760 ;
        RECT  1.880 -0.180 2.220 0.760 ;
        RECT  0.440 -0.180 0.780 1.280 ;
        END
    END VSS
END INV_X32_18_SVT_WB

MACRO INV_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.630 0.985 2.160 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.445 1.540 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  0.440 2.570 0.780 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  0.440 -0.180 0.780 1.230 ;
        END
    END VSS
END INV_X2_18_SVT_WB

MACRO INV_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.356  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.360 1.650 4.475 2.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.996  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.860 2.590 8.200 3.390 ;
        RECT  0.900 0.985 8.200 1.270 ;
        RECT  7.860 0.470 8.200 1.270 ;
        RECT  0.900 2.590 8.200 2.930 ;
        RECT  6.420 2.590 6.760 3.390 ;
        RECT  6.420 0.470 6.760 1.270 ;
        RECT  4.820 0.985 5.720 2.930 ;
        RECT  5.100 0.470 5.440 3.390 ;
        RECT  3.660 2.590 4.000 3.390 ;
        RECT  3.660 0.470 4.000 1.270 ;
        RECT  2.340 2.590 2.680 3.390 ;
        RECT  2.340 0.470 2.680 1.270 ;
        RECT  0.900 2.590 1.240 3.390 ;
        RECT  0.900 0.490 1.240 1.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.140 3.165 7.480 4.100 ;
        RECT  4.380 3.165 4.720 4.100 ;
        RECT  1.620 3.160 1.960 4.100 ;
        RECT  0.180 2.580 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.140 -0.180 7.480 0.755 ;
        RECT  4.380 -0.180 4.720 0.755 ;
        RECT  1.620 -0.180 1.960 0.755 ;
        RECT  0.180 -0.180 0.520 1.280 ;
        END
    END VSS
END INV_X24_18_SVT_WB

MACRO INV_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.715  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.600 2.965 2.170 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.668  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.860 2.570 6.520 2.930 ;
        RECT  0.930 0.950 6.520 1.280 ;
        RECT  4.860 2.570 5.200 3.390 ;
        RECT  4.860 0.470 5.200 1.280 ;
        RECT  0.930 2.570 6.520 2.925 ;
        RECT  3.385 0.950 3.815 2.925 ;
        RECT  2.220 2.570 2.560 3.390 ;
        RECT  2.220 0.470 2.560 1.280 ;
        RECT  0.930 2.570 1.240 3.390 ;
        RECT  0.930 0.470 1.240 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.740 3.565 7.080 4.100 ;
        RECT  2.980 3.560 3.320 4.100 ;
        RECT  0.180 2.580 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.730 -0.180 7.090 0.360 ;
        RECT  2.965 -0.180 3.330 0.360 ;
        RECT  0.180 -0.180 0.520 1.285 ;
        END
    END VSS
END INV_X20_18_SVT_WB

MACRO INV_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.605 1.210 0.985 1.745 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.670 1.540 3.075 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  0.440 2.890 0.780 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  0.440 -0.180 0.780 0.980 ;
        END
    END VSS
END INV_X1_18_SVT_WB

MACRO INV_X18_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X18_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.319  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.625 2.905 2.165 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.346  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.920 2.420 6.540 2.760 ;
        RECT  0.920 0.955 6.540 1.280 ;
        RECT  4.880 2.420 5.220 3.230 ;
        RECT  4.880 0.470 5.220 1.280 ;
        RECT  2.240 2.420 5.220 2.765 ;
        RECT  3.430 0.955 3.820 2.765 ;
        RECT  2.240 2.420 2.580 3.230 ;
        RECT  2.240 0.470 2.580 1.280 ;
        RECT  0.920 0.470 1.275 1.280 ;
        RECT  0.920 2.420 1.260 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  5.635 3.565 5.985 4.100 ;
        RECT  2.995 3.565 3.345 4.100 ;
        RECT  0.200 2.600 0.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  5.640 -0.180 5.980 0.360 ;
        RECT  3.000 -0.180 3.340 0.360 ;
        RECT  0.200 -0.180 0.540 1.330 ;
        END
    END VSS
END INV_X18_18_SVT_WB

MACRO INV_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.046  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.610 2.380 2.205 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.616  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.820 2.450 5.160 3.235 ;
        RECT  0.725 1.050 5.160 1.380 ;
        RECT  4.820 0.470 5.160 1.380 ;
        RECT  0.725 2.450 5.160 2.740 ;
        RECT  3.500 2.450 3.840 3.275 ;
        RECT  3.505 0.555 3.825 1.380 ;
        RECT  2.935 1.050 3.290 2.740 ;
        RECT  2.060 2.450 2.400 3.260 ;
        RECT  2.060 0.470 2.400 1.380 ;
        RECT  0.725 0.900 1.080 1.380 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.540 2.580 5.880 4.100 ;
        RECT  2.780 3.105 3.120 4.100 ;
        RECT  0.180 3.560 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  5.540 -0.180 5.880 1.280 ;
        RECT  2.780 -0.180 3.120 0.780 ;
        RECT  0.180 -0.180 0.520 0.360 ;
        END
    END VSS
END INV_X16_18_SVT_WB

MACRO INV_X14_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X14_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.772  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.625 1.580 2.430 2.200 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.620  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.980 2.475 5.320 3.390 ;
        RECT  0.900 0.995 5.320 1.280 ;
        RECT  4.980 0.470 5.320 1.280 ;
        RECT  0.900 2.475 5.320 2.815 ;
        RECT  3.540 2.475 3.880 3.390 ;
        RECT  3.540 0.470 3.880 1.280 ;
        RECT  0.900 2.475 3.880 2.820 ;
        RECT  2.855 0.995 3.260 2.820 ;
        RECT  2.220 2.475 2.560 3.390 ;
        RECT  2.220 0.470 2.560 1.280 ;
        RECT  0.900 2.475 1.240 3.390 ;
        RECT  0.900 0.470 1.240 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.260 3.075 4.600 4.100 ;
        RECT  0.180 2.580 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.260 -0.180 4.600 0.765 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
END INV_X14_18_SVT_WB

MACRO INV_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.133  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.610 1.620 1.865 2.210 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.294  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.575 3.720 2.945 ;
        RECT  2.365 1.045 3.720 1.385 ;
        RECT  2.365 1.045 2.710 2.945 ;
        RECT  2.060 2.575 2.400 3.390 ;
        RECT  2.060 0.530 2.400 1.380 ;
        RECT  0.740 1.040 2.400 1.380 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.935 3.560 4.290 4.100 ;
        RECT  0.180 3.565 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.930 -0.180 4.295 0.355 ;
        RECT  0.180 -0.180 0.520 0.390 ;
        END
    END VSS
END INV_X12_18_SVT_WB

MACRO INV_X10_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X10_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.600 1.860 2.215 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.317  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.390 2.570 3.730 3.390 ;
        RECT  0.750 0.910 3.730 1.290 ;
        RECT  3.390 0.470 3.730 1.290 ;
        RECT  0.750 2.570 3.730 2.940 ;
        RECT  2.330 0.910 2.690 2.940 ;
        RECT  2.070 0.470 2.415 1.290 ;
        RECT  2.070 2.570 2.410 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.180 3.560 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.180 -0.180 0.505 0.405 ;
        END
    END VSS
END INV_X10_18_SVT_WB

MACRO INV_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.210 0.945 1.590 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.200 0.640 1.545 3.260 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  0.440 2.920 0.780 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  0.440 -0.180 0.780 0.980 ;
        END
    END VSS
END INV_X0_18_SVT_WB

MACRO INV_B_OAI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_OAI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.155 0.860 2.060 ;
        RECT  0.140 1.155 0.860 1.630 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.290 1.475 2.520 ;
        RECT  1.190 1.820 1.475 2.520 ;
        RECT  0.700 2.290 1.080 2.750 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.765 3.325 2.290 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.440 2.630 5.780 3.440 ;
        RECT  4.015 1.155 5.780 1.400 ;
        RECT  5.440 0.485 5.780 1.400 ;
        RECT  4.015 2.630 5.780 2.870 ;
        RECT  4.600 1.155 5.005 2.870 ;
        RECT  4.015 2.630 4.340 3.440 ;
        RECT  4.015 0.515 4.340 1.400 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  6.160 2.630 6.500 4.100 ;
        RECT  4.720 3.100 5.060 4.100 ;
        RECT  3.280 3.110 3.620 4.100 ;
        RECT  0.280 3.110 0.620 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.160 -0.180 6.500 1.280 ;
        RECT  4.720 -0.180 5.060 0.810 ;
        RECT  3.280 -0.180 3.620 0.810 ;
        RECT  1.800 -0.180 2.140 0.405 ;
        RECT  0.280 -0.180 0.620 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.000 0.635 2.250 0.885 ;
        RECT  2.020 0.635 2.250 2.160 ;
        RECT  1.705 1.815 2.250 2.160 ;
        RECT  1.705 1.815 1.935 3.095 ;
        RECT  1.430 2.755 1.935 3.095 ;
        RECT  2.560 0.535 2.900 1.345 ;
        RECT  2.560 1.110 3.785 1.345 ;
        RECT  3.555 1.740 4.100 2.080 ;
        RECT  3.555 1.110 3.785 2.875 ;
        RECT  2.165 2.535 3.785 2.875 ;
        RECT  2.165 2.535 2.470 3.345 ;
    END
END INV_B_OAI21_X8_18_SVT_WB

MACRO INV_B_OAI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_OAI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.460 1.770 0.980 2.210 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.640 1.660 2.055 ;
        RECT  1.210 1.640 1.540 2.150 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.565 3.320 2.100 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.945 2.940 4.915 3.170 ;
        RECT  4.685 0.470 4.915 3.170 ;
        RECT  3.940 0.470 4.915 0.810 ;
        RECT  3.945 2.940 4.390 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.220 3.110 3.560 4.100 ;
        RECT  0.220 2.545 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.220 -0.180 3.560 0.810 ;
        RECT  1.740 -0.180 2.080 0.875 ;
        RECT  0.220 -0.180 0.560 1.345 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.980 0.590 1.320 1.385 ;
        RECT  0.980 1.105 2.270 1.385 ;
        RECT  1.985 1.105 2.270 2.610 ;
        RECT  1.370 2.380 2.270 2.610 ;
        RECT  1.370 2.380 1.710 3.135 ;
        RECT  2.500 0.590 2.840 1.335 ;
        RECT  2.500 1.105 3.930 1.335 ;
        RECT  3.700 1.620 4.455 1.960 ;
        RECT  3.700 1.105 3.930 2.560 ;
        RECT  2.500 2.330 3.930 2.560 ;
        RECT  2.500 2.330 2.730 3.190 ;
        RECT  2.070 2.850 2.730 3.190 ;
    END
END INV_B_OAI21_X4_18_SVT_WB

MACRO INV_B_OAI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_OAI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 2.380 3.445 2.710 ;
        RECT  3.135 1.860 3.445 2.710 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.765 2.905 2.150 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.265 1.820 1.075 2.310 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.920 1.155 2.965 1.440 ;
        RECT  2.195 2.380 2.660 3.385 ;
        RECT  1.920 2.380 2.660 2.630 ;
        RECT  1.920 1.155 2.150 2.630 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.385 3.040 3.725 4.100 ;
        RECT  1.435 3.045 1.775 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.675 -0.180 1.485 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.495 1.080 0.835 1.590 ;
        RECT  0.495 1.360 1.690 1.590 ;
        RECT  1.410 1.360 1.690 2.785 ;
        RECT  0.205 2.555 1.690 2.785 ;
        RECT  0.205 2.555 1.015 3.065 ;
        RECT  1.895 0.610 3.685 0.925 ;
        RECT  3.345 0.610 3.685 1.365 ;
    END
END INV_B_OAI21_X2_18_SVT_WB

MACRO INV_B_OAI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_OAI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.620 3.220 2.430 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.765 1.620 2.200 2.430 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.620 0.700 2.380 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.670 2.890 2.660 3.270 ;
        RECT  2.430 1.050 2.660 3.270 ;
        RECT  2.125 1.050 2.660 1.390 ;
        RECT  1.670 2.660 2.010 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.015 3.515 3.125 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.295 -0.180 1.105 0.595 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 0.995 1.395 1.335 ;
        RECT  1.165 0.995 1.395 2.840 ;
        RECT  0.200 2.610 1.395 2.840 ;
        RECT  0.200 2.610 0.540 2.950 ;
    END
END INV_B_OAI21_X1_18_SVT_WB

MACRO INV_B_OAI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_OAI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.620 3.220 2.430 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.675 2.195 2.430 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.620 0.760 2.380 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.496  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.635 2.660 2.655 3.220 ;
        RECT  2.425 1.100 2.655 3.220 ;
        RECT  2.220 1.100 2.655 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.995 3.450 3.105 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.900 -0.180 1.240 0.900 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.560 0.520 1.365 ;
        RECT  0.180 1.135 1.405 1.365 ;
        RECT  1.120 1.135 1.405 2.840 ;
        RECT  0.180 2.610 1.405 2.840 ;
        RECT  0.180 2.610 0.520 2.950 ;
    END
END INV_B_OAI21_X0_18_SVT_WB

MACRO INV_B_AOI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_AOI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.290 0.860 2.765 ;
        RECT  0.520 1.860 0.860 2.765 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.190 1.400 1.475 1.960 ;
        RECT  0.700 1.400 1.475 1.630 ;
        RECT  0.700 1.170 1.080 1.630 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.620 3.325 2.100 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.440 2.420 5.780 3.230 ;
        RECT  4.015 1.050 5.780 1.290 ;
        RECT  5.440 0.480 5.780 1.290 ;
        RECT  4.015 2.420 5.780 2.765 ;
        RECT  4.600 1.050 5.005 2.765 ;
        RECT  4.015 2.420 4.340 3.230 ;
        RECT  4.015 0.480 4.340 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  6.160 2.640 6.500 4.100 ;
        RECT  4.720 3.110 5.060 4.100 ;
        RECT  3.280 3.110 3.620 4.100 ;
        RECT  1.800 3.515 2.140 4.100 ;
        RECT  0.280 3.110 0.620 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.160 -0.180 6.500 1.290 ;
        RECT  4.720 -0.180 5.060 0.820 ;
        RECT  3.280 -0.180 3.620 0.810 ;
        RECT  0.280 -0.180 0.620 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.430 0.825 1.935 1.165 ;
        RECT  1.705 0.825 1.935 1.965 ;
        RECT  1.705 1.620 2.250 1.965 ;
        RECT  2.020 1.620 2.250 3.285 ;
        RECT  1.000 3.035 2.250 3.285 ;
        RECT  2.165 0.575 2.470 1.385 ;
        RECT  2.165 1.045 3.785 1.385 ;
        RECT  3.555 1.840 4.100 2.180 ;
        RECT  3.555 1.045 3.785 2.810 ;
        RECT  2.560 2.575 3.785 2.810 ;
        RECT  2.560 2.575 2.900 3.385 ;
    END
END INV_B_AOI21_X8_18_SVT_WB

MACRO INV_B_AOI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_AOI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.620 0.935 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.165 2.295 1.715 2.710 ;
        RECT  1.165 1.840 1.495 2.710 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.895 1.615 3.280 2.150 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 2.920 4.805 3.385 ;
        RECT  4.575 0.500 4.805 3.385 ;
        RECT  3.895 0.500 4.805 0.805 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.180 3.090 3.580 4.100 ;
        RECT  1.700 3.515 2.040 4.100 ;
        RECT  0.180 2.565 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.180 -0.180 3.580 0.775 ;
        RECT  0.180 -0.180 0.520 1.390 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.330 0.630 1.670 1.610 ;
        RECT  1.330 1.380 2.230 1.610 ;
        RECT  1.945 1.380 2.230 3.285 ;
        RECT  0.900 3.035 2.230 3.285 ;
        RECT  2.030 0.475 2.690 0.815 ;
        RECT  2.460 0.475 2.690 1.385 ;
        RECT  2.460 1.045 4.040 1.385 ;
        RECT  3.780 1.045 4.040 2.685 ;
        RECT  2.460 2.380 4.040 2.685 ;
        RECT  2.460 2.380 2.800 3.385 ;
    END
END INV_B_AOI21_X4_18_SVT_WB

MACRO INV_B_AOI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_AOI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.985 1.260 3.270 1.960 ;
        RECT  2.755 1.260 3.270 1.590 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 1.820 2.755 2.205 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.585 1.260 1.030 1.725 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.435 2.725 2.775 ;
        RECT  1.955 0.535 2.295 1.540 ;
        RECT  1.770 0.830 2.000 2.775 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.905 3.515 1.245 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.105 -0.180 3.445 0.810 ;
        RECT  1.195 -0.180 1.535 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.435 0.690 1.540 1.030 ;
        RECT  1.260 0.690 1.540 2.720 ;
        RECT  0.345 2.380 1.540 2.720 ;
        RECT  3.105 2.435 3.445 3.255 ;
        RECT  1.655 3.015 3.445 3.255 ;
    END
END INV_B_AOI21_X2_18_SVT_WB

MACRO INV_B_AOI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_AOI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.910 1.495 3.220 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.715 1.680 2.150 2.145 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.475 1.625 0.980 2.235 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.155 2.455 2.660 2.795 ;
        RECT  2.380 0.900 2.660 2.795 ;
        RECT  1.710 0.900 2.660 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.795 3.515 1.135 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.020 -0.180 3.160 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.235 1.055 1.480 1.395 ;
        RECT  1.250 1.055 1.480 3.095 ;
        RECT  0.235 2.755 1.480 3.095 ;
    END
END INV_B_AOI21_X1_18_SVT_WB

MACRO INV_B_AOI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_B_AOI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 1.210 3.235 1.810 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.565 2.150 2.100 ;
        END
    END A1
    PIN B0N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.525 0.505 2.150 ;
        END
    END B0N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 2.380 2.710 2.720 ;
        RECT  2.380 0.950 2.610 2.720 ;
        RECT  1.660 0.950 2.610 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.900 3.050 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.940 -0.180 3.170 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.950 1.430 1.290 ;
        RECT  1.090 0.950 1.430 2.815 ;
        RECT  0.180 2.475 1.430 2.815 ;
        RECT  0.180 2.475 0.520 3.390 ;
    END
END INV_B_AOI21_X0_18_SVT_WB

MACRO INV_A_OAI22_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI22_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.255 2.880 2.770 3.220 ;
        RECT  2.255 1.775 2.540 3.220 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.475 1.665 5.425 2.160 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.210 1.515 2.080 ;
        RECT  0.615 1.210 1.515 1.620 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.285 0.890 2.520 ;
        RECT  0.550 1.850 0.890 2.520 ;
        RECT  0.140 2.285 0.540 2.775 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.775 2.545 11.115 3.385 ;
        RECT  9.225 1.055 11.115 1.350 ;
        RECT  10.775 0.535 11.115 1.350 ;
        RECT  9.225 2.545 11.115 2.940 ;
        RECT  10.130 1.055 10.530 2.940 ;
        RECT  9.225 0.590 9.575 1.350 ;
        RECT  9.225 2.545 9.565 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.495 2.545 11.830 4.100 ;
        RECT  9.980 3.560 10.365 4.100 ;
        RECT  8.460 3.570 8.800 4.100 ;
        RECT  4.040 3.095 4.380 4.100 ;
        RECT  3.140 3.110 3.480 4.100 ;
        RECT  0.310 3.110 0.650 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.500 -0.180 11.870 1.360 ;
        RECT  9.990 -0.180 10.360 0.360 ;
        RECT  8.460 -0.180 8.800 0.350 ;
        RECT  3.910 -0.180 4.250 0.350 ;
        RECT  0.940 -0.180 1.280 0.355 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.595 3.480 0.825 ;
        RECT  4.760 1.085 6.420 1.390 ;
        RECT  2.890 1.860 3.270 2.660 ;
        RECT  5.655 1.085 6.020 2.920 ;
        RECT  2.890 2.400 4.205 2.660 ;
        RECT  3.950 2.570 6.420 2.845 ;
        RECT  4.760 2.570 6.420 2.920 ;
        RECT  4.760 2.570 5.100 3.390 ;
        RECT  6.080 2.570 6.420 3.390 ;
        RECT  3.810 0.580 7.580 0.810 ;
        RECT  3.810 0.580 4.040 1.345 ;
        RECT  1.750 1.105 4.040 1.345 ;
        RECT  7.285 0.580 7.580 2.050 ;
        RECT  7.285 1.750 8.020 2.050 ;
        RECT  1.750 1.105 2.025 3.295 ;
        RECT  7.900 0.905 8.585 1.160 ;
        RECT  8.250 0.905 8.585 2.670 ;
        RECT  8.250 1.620 9.765 1.960 ;
        RECT  8.250 1.620 8.590 2.670 ;
        RECT  7.900 2.405 8.590 2.670 ;
    END
END INV_A_OAI22_X8_18_SVT_WB

MACRO INV_A_OAI22_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI22_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.670 3.365 2.150 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.820 1.195 2.355 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.770 1.200 6.580 1.905 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.105 2.135 7.275 2.365 ;
        RECT  6.910 1.860 7.275 2.365 ;
        RECT  5.105 1.620 5.460 2.365 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.760 2.890 6.340 3.295 ;
        RECT  4.645 2.595 6.340 3.295 ;
        RECT  4.645 1.100 4.875 3.295 ;
        RECT  2.355 1.100 4.875 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  7.150 2.695 7.505 4.100 ;
        RECT  4.410 3.525 4.750 4.100 ;
        RECT  1.600 3.160 1.940 4.100 ;
        RECT  0.165 2.685 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.240 -0.180 5.580 0.350 ;
        RECT  0.180 -0.180 0.520 1.355 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.610 1.240 1.590 ;
        RECT  0.900 1.360 2.125 1.590 ;
        RECT  1.855 2.380 4.415 2.610 ;
        RECT  3.900 2.150 4.415 2.610 ;
        RECT  4.130 1.840 4.415 2.610 ;
        RECT  1.855 1.360 2.125 2.875 ;
        RECT  0.900 2.610 2.125 2.875 ;
        RECT  0.900 2.610 1.240 3.385 ;
        RECT  1.600 0.580 7.660 0.870 ;
        RECT  7.320 0.580 7.660 1.345 ;
    END
END INV_A_OAI22_X4_18_SVT_WB

MACRO INV_A_OAI22_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI22_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.295 1.745 2.710 2.290 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.535 0.560 2.155 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.510 3.305 2.235 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.765 1.665 4.340 2.205 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.916  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.605 2.880 3.105 3.220 ;
        RECT  1.805 1.100 2.395 1.435 ;
        RECT  1.805 1.100 2.060 3.220 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.925 2.435 4.265 4.100 ;
        RECT  0.235 3.570 1.640 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.395 -0.180 3.735 1.280 ;
        RECT  0.235 -0.180 0.575 0.375 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.850 1.740 1.575 2.160 ;
        RECT  0.850 0.965 1.080 2.720 ;
    END
END INV_A_OAI22_X2_18_SVT_WB

MACRO INV_A_OAI22_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI22_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.665 2.660 2.410 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.210 0.510 2.020 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 2.375 3.675 2.750 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.005 1.620 4.340 2.285 ;
        RECT  3.650 1.620 4.340 1.975 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.540 2.980 2.940 3.285 ;
        RECT  1.885 1.045 2.350 1.385 ;
        RECT  1.540 2.915 2.275 3.285 ;
        RECT  1.885 1.045 2.115 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.750 2.985 4.090 4.100 ;
        RECT  0.180 3.570 1.590 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.320 -0.180 3.660 1.335 ;
        RECT  0.175 -0.180 0.525 0.355 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.875 1.070 2.430 ;
        RECT  0.740 2.080 1.655 2.430 ;
        RECT  0.740 0.875 1.065 2.965 ;
    END
END INV_A_OAI22_X1_18_SVT_WB

MACRO INV_A_OAI22_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI22_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.335 1.615 2.690 2.440 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.640 0.520 2.210 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.560 3.410 2.190 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.835 1.770 4.340 2.420 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.580  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.830 2.785 3.285 3.220 ;
        RECT  1.875 1.040 2.360 1.375 ;
        RECT  1.875 1.040 2.105 3.220 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.890 3.570 4.230 4.100 ;
        RECT  1.440 3.570 1.780 4.100 ;
        RECT  0.180 3.565 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.330 -0.180 3.670 1.330 ;
        RECT  0.180 -0.180 0.520 0.365 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.750 0.990 1.080 2.200 ;
        RECT  0.750 1.855 1.645 2.200 ;
        RECT  0.750 0.990 1.075 3.120 ;
    END
END INV_A_OAI22_X0_18_SVT_WB

MACRO INV_A_OAI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.960 2.700 2.710 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.189  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.255 0.500 2.820 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.378  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.765 1.670 2.300 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.305 2.545 7.645 3.385 ;
        RECT  5.985 1.055 7.645 1.350 ;
        RECT  7.305 0.535 7.645 1.350 ;
        RECT  5.985 2.545 7.645 2.940 ;
        RECT  6.780 1.055 7.155 2.940 ;
        RECT  5.985 0.590 6.335 1.350 ;
        RECT  5.985 2.545 6.325 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  5.220 3.570 5.560 4.100 ;
        RECT  3.390 2.530 3.675 4.100 ;
        RECT  1.105 3.515 1.445 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  5.220 -0.180 5.560 0.350 ;
        RECT  1.105 -0.180 1.445 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.340 1.065 0.960 1.405 ;
        RECT  2.930 1.960 3.405 2.300 ;
        RECT  0.730 1.065 0.960 3.280 ;
        RECT  2.930 1.960 3.160 3.280 ;
        RECT  0.345 3.050 3.160 3.280 ;
        RECT  0.345 3.050 0.685 3.385 ;
        RECT  1.830 0.535 3.655 0.785 ;
        RECT  1.900 1.085 4.350 1.340 ;
        RECT  4.045 1.085 4.350 2.090 ;
        RECT  4.045 1.750 4.780 2.090 ;
        RECT  1.900 1.085 2.150 2.820 ;
        RECT  4.660 0.905 5.345 1.160 ;
        RECT  5.010 0.905 5.345 2.670 ;
        RECT  5.010 1.620 6.525 1.960 ;
        RECT  5.010 1.620 5.350 2.670 ;
        RECT  4.660 2.405 5.350 2.670 ;
    END
END INV_A_OAI21_X8_18_SVT_WB

MACRO INV_A_OAI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.630 2.180 2.175 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.207  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.770 0.495 2.445 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.205 1.595 1.540 2.200 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.080 2.585 6.020 2.910 ;
        RECT  5.695 1.050 6.020 2.910 ;
        RECT  5.080 1.050 6.020 1.345 ;
        RECT  5.080 2.585 5.430 3.385 ;
        RECT  5.080 0.535 5.415 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.320 3.515 4.660 4.100 ;
        RECT  3.100 3.565 3.440 4.100 ;
        RECT  0.860 3.515 1.200 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.320 -0.180 4.660 0.350 ;
        RECT  0.860 -0.180 1.200 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 1.155 0.960 1.540 ;
        RECT  0.180 2.675 0.960 2.910 ;
        RECT  0.730 1.155 0.960 3.280 ;
        RECT  2.870 1.860 3.160 3.280 ;
        RECT  0.730 3.050 3.160 3.280 ;
        RECT  1.620 0.470 3.400 0.755 ;
        RECT  2.335 0.985 3.530 1.220 ;
        RECT  3.300 0.985 3.530 1.630 ;
        RECT  3.300 1.325 4.145 1.630 ;
        RECT  3.815 1.325 4.145 2.180 ;
        RECT  3.815 1.865 4.390 2.180 ;
        RECT  2.410 0.985 2.640 2.820 ;
        RECT  1.675 2.470 2.640 2.820 ;
        RECT  3.760 0.800 4.850 1.095 ;
        RECT  4.620 1.615 5.265 2.000 ;
        RECT  4.620 0.800 4.850 2.750 ;
        RECT  3.760 2.410 4.850 2.750 ;
    END
END INV_A_OAI21_X4_18_SVT_WB

MACRO INV_A_OAI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.860 2.700 2.710 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.990 0.500 2.790 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.765 1.670 2.345 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.900 1.155 3.305 1.540 ;
        RECT  1.900 1.155 2.150 2.820 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.390 2.530 3.675 4.100 ;
        RECT  1.105 3.515 1.445 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.105 -0.180 1.445 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.340 1.075 0.960 1.415 ;
        RECT  2.930 1.860 3.405 2.200 ;
        RECT  0.730 1.075 0.960 3.280 ;
        RECT  2.930 1.860 3.160 3.280 ;
        RECT  0.345 3.050 3.160 3.280 ;
        RECT  0.345 3.050 0.685 3.385 ;
        RECT  1.865 0.535 3.645 0.875 ;
    END
END INV_A_OAI21_X2_18_SVT_WB

MACRO INV_A_OAI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.650 2.130 2.460 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.770 0.980 2.325 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.230 1.580 2.660 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 2.940 2.770 3.285 ;
        RECT  2.360 2.935 2.770 3.285 ;
        RECT  2.360 1.060 2.590 3.285 ;
        RECT  2.200 1.060 2.590 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.000 2.975 1.340 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.840 -0.180 1.180 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.580 3.160 0.810 ;
        RECT  0.115 0.580 0.620 1.365 ;
        RECT  2.820 0.580 3.160 2.040 ;
        RECT  0.115 0.580 0.345 3.285 ;
        RECT  0.115 2.945 0.620 3.285 ;
    END
END INV_A_OAI21_X1_18_SVT_WB

MACRO INV_A_OAI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.795 1.760 2.150 2.330 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.820 1.070 2.100 ;
        RECT  0.575 1.820 0.860 2.490 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.185 2.315 1.565 2.850 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 3.045 2.660 3.385 ;
        RECT  2.380 1.080 2.660 3.385 ;
        RECT  2.200 1.080 2.660 1.410 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.000 3.080 1.340 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.840 -0.180 1.180 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.605 3.195 0.835 ;
        RECT  0.115 0.605 0.620 1.145 ;
        RECT  2.890 0.605 3.195 2.060 ;
        RECT  0.115 0.605 0.345 3.385 ;
        RECT  0.115 3.045 0.620 3.385 ;
    END
END INV_A_OAI21_X0_18_SVT_WB

MACRO INV_A_OAI211_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI211_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.695 1.420 4.340 1.680 ;
        RECT  4.060 1.200 4.340 1.680 ;
        RECT  3.695 1.420 3.940 1.960 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.465 1.770 0.980 2.200 ;
        RECT  0.465 1.390 0.810 2.200 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.620 2.320 2.210 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.260 1.590 1.600 ;
        RECT  1.230 1.260 1.515 1.960 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.180 0.535 6.615 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.420 3.515 5.760 4.100 ;
        RECT  2.445 3.555 2.815 4.100 ;
        RECT  0.400 3.460 1.210 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  5.420 -0.180 5.760 0.875 ;
        RECT  1.050 -0.180 1.390 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.310 0.765 2.050 1.030 ;
        RECT  1.820 0.765 2.050 1.390 ;
        RECT  0.310 0.765 0.650 1.105 ;
        RECT  1.820 1.105 2.780 1.390 ;
        RECT  2.550 1.840 3.005 2.180 ;
        RECT  2.550 1.105 2.780 2.710 ;
        RECT  0.310 2.440 2.780 2.710 ;
        RECT  0.310 2.440 0.650 2.780 ;
        RECT  2.280 0.520 2.580 0.860 ;
        RECT  2.280 0.630 4.020 0.860 ;
        RECT  3.680 0.630 4.020 0.970 ;
        RECT  3.010 1.100 3.465 1.440 ;
        RECT  4.870 1.885 5.240 2.180 ;
        RECT  4.255 1.950 5.240 2.180 ;
        RECT  3.235 1.100 3.465 3.280 ;
        RECT  4.255 1.950 4.485 2.760 ;
        RECT  3.235 2.525 4.485 2.760 ;
        RECT  3.235 2.525 4.020 3.280 ;
        RECT  1.700 2.940 4.020 3.280 ;
        RECT  4.660 0.535 5.000 1.485 ;
        RECT  4.660 1.255 5.950 1.485 ;
        RECT  5.720 1.255 5.950 2.750 ;
        RECT  4.715 2.410 5.950 2.750 ;
        RECT  4.715 2.410 5.000 3.385 ;
    END
END INV_A_OAI211_X4_18_SVT_WB

MACRO INV_A_OAI211_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI211_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.695 1.420 4.340 1.680 ;
        RECT  4.060 1.200 4.340 1.680 ;
        RECT  3.695 1.420 3.940 1.960 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.465 1.770 0.980 2.200 ;
        RECT  0.465 1.390 0.810 2.200 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.620 2.320 2.210 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.260 1.590 1.600 ;
        RECT  1.230 1.260 1.515 1.960 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.821  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 2.940 4.020 3.280 ;
        RECT  3.235 2.525 4.020 3.280 ;
        RECT  3.235 1.100 3.465 3.280 ;
        RECT  3.010 1.100 3.465 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  2.445 3.555 2.815 4.100 ;
        RECT  0.400 3.460 1.210 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  1.050 -0.180 1.390 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.310 0.765 2.050 1.030 ;
        RECT  1.820 0.765 2.050 1.390 ;
        RECT  0.310 0.765 0.650 1.105 ;
        RECT  1.820 1.105 2.780 1.390 ;
        RECT  2.550 1.840 3.005 2.180 ;
        RECT  2.550 1.105 2.780 2.710 ;
        RECT  0.310 2.440 2.780 2.710 ;
        RECT  0.310 2.440 0.650 2.780 ;
        RECT  2.280 0.520 2.580 0.860 ;
        RECT  2.280 0.630 4.020 0.860 ;
        RECT  3.680 0.630 4.020 0.970 ;
    END
END INV_A_OAI211_X2_18_SVT_WB

MACRO INV_A_OAI211_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI211_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.760 3.830 2.335 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 1.095 1.030 1.540 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.130 2.230 1.570 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.095 1.540 1.820 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.915  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.865 2.890 4.340 3.360 ;
        RECT  1.565 2.995 4.340 3.225 ;
        RECT  2.990 2.890 4.340 3.225 ;
        RECT  2.990 1.060 3.255 1.400 ;
        RECT  2.990 1.060 3.220 3.225 ;
        RECT  1.565 2.995 1.850 3.275 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  2.325 3.570 2.665 4.100 ;
        RECT  0.805 3.570 1.145 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  0.995 -0.180 1.225 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.630 0.520 0.865 ;
        RECT  0.180 0.635 2.760 0.865 ;
        RECT  2.530 0.635 2.760 2.760 ;
        RECT  0.300 2.530 2.760 2.760 ;
        RECT  0.300 2.530 0.530 3.115 ;
    END
END INV_A_OAI211_X1_18_SVT_WB

MACRO INV_A_OAI211_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_OAI211_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.385 1.620 3.780 2.390 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.460 0.745 1.880 ;
        RECT  0.140 1.460 0.510 2.215 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.590 1.105 2.130 1.590 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.820 1.625 2.245 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.500 3.050 3.710 3.280 ;
        RECT  2.925 2.620 3.710 3.280 ;
        RECT  2.925 1.100 3.155 3.280 ;
        RECT  2.870 1.100 3.155 1.440 ;
        RECT  1.500 3.050 1.840 3.380 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  2.260 3.510 3.070 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.740 -0.180 1.080 0.415 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.645 2.640 0.875 ;
        RECT  0.180 0.645 0.520 1.205 ;
        RECT  2.410 0.645 2.640 2.820 ;
        RECT  2.410 1.905 2.695 2.820 ;
        RECT  0.180 2.590 2.695 2.820 ;
        RECT  0.180 2.590 0.520 3.380 ;
    END
END INV_A_OAI211_X0_18_SVT_WB

MACRO INV_A_NOR4_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR4_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.640 2.150 1.030 2.745 ;
        RECT  0.640 1.790 0.925 2.745 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 1.820 5.240 2.280 ;
        RECT  4.190 1.455 4.530 2.280 ;
        RECT  2.900 1.455 4.530 1.685 ;
        RECT  2.900 1.455 3.240 2.005 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.610 0.995 5.950 2.060 ;
        RECT  5.130 0.995 5.950 1.555 ;
        RECT  2.230 0.995 5.950 1.225 ;
        RECT  2.230 0.995 2.570 2.005 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 2.695 6.705 2.925 ;
        RECT  6.400 1.830 6.705 2.925 ;
        RECT  1.260 1.810 1.540 2.925 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.186  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.940 3.155 7.165 3.450 ;
        RECT  6.935 1.200 7.165 3.450 ;
        RECT  6.180 1.200 7.165 1.540 ;
        RECT  6.180 0.510 6.520 1.540 ;
        RECT  1.620 0.510 6.520 0.765 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  1.065 3.155 1.405 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  0.900 -0.180 1.240 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.570 0.520 1.500 ;
        RECT  0.180 1.160 2.000 1.500 ;
        RECT  1.770 1.160 2.000 2.465 ;
        RECT  3.620 1.915 3.960 2.465 ;
        RECT  1.770 2.235 3.960 2.465 ;
        RECT  0.180 0.570 0.410 3.450 ;
        RECT  0.180 3.110 0.685 3.450 ;
    END
END INV_A_NOR4_X4_18_SVT_WB

MACRO INV_A_NOR4_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR4_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.595 1.695 1.030 2.275 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.710 1.725 3.220 2.295 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.720 2.305 2.195 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.705 1.590 2.515 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.939  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.915 0.640 4.200 3.290 ;
        RECT  1.680 0.640 4.200 0.980 ;
        RECT  3.200 0.535 3.540 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  0.990 3.515 1.330 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.960 -0.180 4.300 0.405 ;
        RECT  2.440 -0.180 2.780 0.405 ;
        RECT  0.920 -0.180 1.260 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.360 1.040 0.720 1.440 ;
        RECT  0.360 1.210 3.685 1.440 ;
        RECT  0.360 2.550 0.700 3.120 ;
        RECT  3.450 1.210 3.685 3.120 ;
        RECT  0.360 2.890 3.685 3.120 ;
    END
END INV_A_NOR4_X2_18_SVT_WB

MACRO INV_A_NOR4_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR4_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.115 0.480 2.710 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.225 2.330 2.660 2.795 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.570 2.240 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 2.480 1.790 2.710 ;
        RECT  1.220 2.200 1.560 2.710 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.873  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.350 2.890 3.805 3.270 ;
        RECT  3.575 0.950 3.805 3.270 ;
        RECT  1.520 0.950 3.805 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.050 -0.180 3.675 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 0.990 1.440 ;
        RECT  2.890 2.190 3.345 2.530 ;
        RECT  0.710 1.100 0.990 3.270 ;
        RECT  0.180 2.940 0.990 3.270 ;
        RECT  2.890 2.190 3.120 3.270 ;
        RECT  0.180 3.040 3.120 3.270 ;
    END
END INV_A_NOR4_X1_18_SVT_WB

MACRO INV_A_NOR4_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR4_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.980 0.760 2.740 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.260 2.330 2.695 2.795 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.785 2.390 2.100 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.205 2.300 1.610 2.800 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.385 2.890 3.785 3.310 ;
        RECT  3.555 0.805 3.785 3.310 ;
        RECT  1.500 0.805 3.785 1.095 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.030 3.540 1.370 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.860 -0.180 3.740 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.805 0.520 1.555 ;
        RECT  0.180 1.325 3.325 1.555 ;
        RECT  2.925 1.325 3.325 2.135 ;
        RECT  0.180 2.970 0.520 3.310 ;
        RECT  2.925 1.325 3.155 3.310 ;
        RECT  0.180 3.030 3.155 3.310 ;
    END
END INV_A_NOR4_X0_18_SVT_WB

MACRO INV_A_NOR3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.695 1.625 1.080 2.150 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.920 1.455 4.340 2.150 ;
        RECT  2.100 1.455 4.340 1.685 ;
        RECT  2.100 1.455 2.440 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.620 0.995 4.960 1.960 ;
        RECT  1.455 0.995 4.960 1.225 ;
        RECT  1.455 0.995 1.740 1.960 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.322  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.010 2.925 5.420 3.265 ;
        RECT  5.190 0.470 5.420 3.265 ;
        RECT  1.620 0.470 5.420 0.765 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.870 3.495 5.210 4.100 ;
        RECT  1.150 3.045 1.490 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  0.895 -0.180 1.225 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.525 0.520 1.280 ;
        RECT  0.180 0.525 0.465 3.190 ;
        RECT  2.770 1.915 3.580 2.695 ;
        RECT  0.180 2.380 3.580 2.695 ;
        RECT  0.180 2.380 0.730 3.190 ;
    END
END INV_A_NOR3_X4_18_SVT_WB

MACRO INV_A_NOR3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.585 2.100 2.200 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.645 1.540 2.200 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.623  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.790 2.480 3.240 3.370 ;
        RECT  3.010 0.535 3.240 3.370 ;
        RECT  2.840 0.535 3.240 1.510 ;
        RECT  1.500 0.535 3.240 0.885 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.820 3.515 1.160 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.115 2.560 1.355 ;
        RECT  2.330 1.740 2.780 2.080 ;
        RECT  2.330 1.115 2.560 2.880 ;
        RECT  0.180 2.540 2.560 2.880 ;
    END
END INV_A_NOR3_X2_18_SVT_WB

MACRO INV_A_NOR3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.730 0.930 2.505 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.730 2.165 2.245 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.165 2.185 1.540 2.725 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.892  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.855 3.060 3.195 3.400 ;
        RECT  2.965 0.700 3.195 3.400 ;
        RECT  1.510 0.700 3.195 1.040 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.940 3.475 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.280 -0.180 1.090 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.810 0.520 1.500 ;
        RECT  0.180 1.270 2.735 1.500 ;
        RECT  2.395 1.270 2.735 2.140 ;
        RECT  0.180 2.905 0.520 3.245 ;
        RECT  2.395 1.270 2.625 3.245 ;
        RECT  0.180 2.955 2.625 3.245 ;
    END
END INV_A_NOR3_X1_18_SVT_WB

MACRO INV_A_NOR3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.340 1.755 0.680 2.565 ;
        RECT  0.140 1.755 0.680 2.150 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.475 2.535 2.105 2.810 ;
        RECT  1.820 1.785 2.105 2.810 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.820 1.590 2.305 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.689  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.795 2.775 3.225 3.115 ;
        RECT  2.995 0.700 3.225 3.115 ;
        RECT  1.510 0.700 3.225 1.095 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.810 3.515 1.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.940 -0.180 1.750 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.805 0.520 1.315 ;
        RECT  0.180 1.085 1.175 1.315 ;
        RECT  0.835 1.085 1.175 1.555 ;
        RECT  0.835 1.325 2.765 1.555 ;
        RECT  2.335 1.325 2.765 2.135 ;
        RECT  0.180 2.795 0.520 3.270 ;
        RECT  2.335 1.325 2.565 3.270 ;
        RECT  0.180 3.040 2.565 3.270 ;
    END
END INV_A_NOR3_X0_18_SVT_WB

MACRO INV_A_NOR2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.790 0.600 2.760 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.220 1.455 6.700 2.120 ;
        RECT  1.840 1.455 6.700 1.685 ;
        RECT  3.980 1.455 4.320 2.005 ;
        RECT  1.840 1.455 2.180 2.005 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.510  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.780 2.695 7.165 2.925 ;
        RECT  6.930 0.985 7.165 2.925 ;
        RECT  2.040 0.995 7.165 1.225 ;
        RECT  3.460 0.985 7.165 1.225 ;
        RECT  6.115 0.495 6.505 1.225 ;
        RECT  5.420 2.695 5.760 3.450 ;
        RECT  4.775 0.470 5.210 1.225 ;
        RECT  3.460 0.455 3.880 1.225 ;
        RECT  2.780 2.695 3.120 3.405 ;
        RECT  2.040 0.485 2.430 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.760 3.155 7.100 4.100 ;
        RECT  4.220 3.155 4.560 4.100 ;
        RECT  1.630 3.110 1.970 4.100 ;
        RECT  0.190 3.110 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  2.745 -0.180 3.170 0.765 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.585 1.250 1.395 ;
        RECT  2.540 1.915 2.880 2.465 ;
        RECT  5.200 1.915 5.540 2.465 ;
        RECT  0.910 2.235 5.540 2.465 ;
        RECT  0.910 0.585 1.250 3.450 ;
    END
END INV_A_NOR2_X8_18_SVT_WB

MACRO INV_A_NOR2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.515 0.570 2.150 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.880 1.455 3.345 2.125 ;
        RECT  1.260 1.455 3.345 1.685 ;
        RECT  1.260 1.455 1.600 1.960 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.755  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.150 2.845 3.805 3.450 ;
        RECT  3.575 0.885 3.805 3.450 ;
        RECT  1.500 0.885 3.805 1.225 ;
        RECT  2.820 0.470 3.160 1.225 ;
        RECT  1.500 0.475 1.840 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.940 3.015 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.270 -0.180 1.080 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.995 1.030 1.285 ;
        RECT  0.800 0.995 1.030 2.615 ;
        RECT  1.980 1.915 2.320 2.615 ;
        RECT  0.180 2.385 2.320 2.615 ;
        RECT  0.180 2.385 0.575 3.455 ;
    END
END INV_A_NOR2_X4_18_SVT_WB

MACRO INV_A_NOR2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.330 0.980 2.710 ;
        RECT  0.700 1.670 0.930 2.710 ;
        RECT  0.355 1.670 0.930 2.010 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.710 1.590 2.180 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.383  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.640 2.585 3.330 ;
        RECT  1.515 0.640 2.585 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.410 3.460 1.110 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.275 -0.180 2.615 0.410 ;
        RECT  0.285 -0.180 1.095 0.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.195 1.100 0.535 1.440 ;
        RECT  0.195 1.210 2.060 1.440 ;
        RECT  0.185 2.380 0.470 3.170 ;
        RECT  1.820 1.210 2.060 3.170 ;
        RECT  0.185 2.940 2.060 3.170 ;
    END
END INV_A_NOR2_X2_18_SVT_WB

MACRO INV_A_NOR2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.685 0.760 2.410 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.195 1.820 1.605 2.410 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.559  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.295 0.700 2.525 3.160 ;
        RECT  1.520 0.700 2.525 0.995 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  1.050 3.100 1.390 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.280 -0.180 2.620 0.460 ;
        RECT  0.290 -0.180 1.100 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.810 0.520 1.455 ;
        RECT  0.180 1.225 2.065 1.455 ;
        RECT  1.785 1.225 2.065 1.670 ;
        RECT  1.835 1.225 2.065 2.870 ;
        RECT  0.290 2.640 2.065 2.870 ;
        RECT  0.290 2.640 0.630 3.005 ;
    END
END INV_A_NOR2_X1_18_SVT_WB

MACRO INV_A_NOR2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.470 0.670 2.300 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.585 1.455 9.965 2.175 ;
        RECT  2.000 1.455 9.965 1.685 ;
        RECT  7.020 1.455 7.360 2.005 ;
        RECT  4.620 1.455 4.960 2.005 ;
        RECT  2.000 1.455 2.340 2.005 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.265  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.195 0.940 10.500 2.870 ;
        RECT  8.680 2.500 10.500 2.870 ;
        RECT  2.220 0.995 10.500 1.225 ;
        RECT  7.980 0.940 10.500 1.225 ;
        RECT  9.400 0.465 9.740 1.225 ;
        RECT  8.680 2.500 9.020 3.310 ;
        RECT  2.940 2.695 9.020 2.935 ;
        RECT  7.980 0.470 8.320 1.225 ;
        RECT  5.100 0.990 10.500 1.225 ;
        RECT  6.540 0.470 6.880 1.225 ;
        RECT  5.100 0.470 5.440 1.225 ;
        RECT  2.220 0.940 4.000 1.225 ;
        RECT  3.660 0.470 4.000 1.225 ;
        RECT  2.940 2.695 3.290 3.450 ;
        RECT  2.220 0.470 2.560 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  10.120 3.110 10.460 4.100 ;
        RECT  7.260 3.165 7.600 4.100 ;
        RECT  4.380 3.165 4.720 4.100 ;
        RECT  1.620 3.110 1.960 4.100 ;
        RECT  0.180 3.110 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  7.260 -0.180 7.600 0.760 ;
        RECT  5.820 -0.180 6.160 0.760 ;
        RECT  4.380 -0.180 4.720 0.760 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  8.045 1.915 8.685 2.200 ;
        RECT  2.700 1.915 3.040 2.465 ;
        RECT  5.600 1.915 5.940 2.465 ;
        RECT  8.045 1.915 8.425 2.465 ;
        RECT  0.900 2.235 8.425 2.465 ;
        RECT  0.900 0.470 1.240 3.450 ;
    END
END INV_A_NOR2_X12_18_SVT_WB

MACRO INV_A_NOR2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NOR2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.600 0.760 2.150 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 2.380 1.605 2.825 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.295 1.140 2.660 3.380 ;
        RECT  1.520 1.140 2.660 1.370 ;
        RECT  1.520 0.860 1.860 1.370 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  1.050 3.515 1.390 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.280 -0.180 2.620 0.820 ;
        RECT  0.760 -0.180 1.100 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.860 0.520 1.370 ;
        RECT  0.180 1.140 1.290 1.370 ;
        RECT  0.990 1.140 1.290 1.830 ;
        RECT  0.990 1.600 2.065 1.830 ;
        RECT  1.750 1.600 2.065 2.110 ;
        RECT  1.835 1.600 2.065 3.285 ;
        RECT  0.290 3.055 2.065 3.285 ;
        RECT  0.290 3.055 0.630 3.380 ;
    END
END INV_A_NOR2_X0_18_SVT_WB

MACRO INV_A_NAND4_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND4_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.640 1.260 1.030 1.600 ;
        RECT  0.640 1.260 0.925 1.960 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.190 1.640 5.240 2.100 ;
        RECT  2.900 2.135 4.530 2.365 ;
        RECT  4.190 1.640 4.530 2.365 ;
        RECT  2.900 1.915 3.240 2.365 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 2.595 5.950 2.825 ;
        RECT  5.610 1.860 5.950 2.825 ;
        RECT  5.130 2.365 5.950 2.825 ;
        RECT  2.230 1.915 2.570 2.825 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.400 0.995 6.705 1.980 ;
        RECT  1.260 0.995 6.705 1.225 ;
        RECT  1.260 0.995 1.540 1.960 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.135  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.180 2.380 7.165 2.720 ;
        RECT  6.935 0.470 7.165 2.720 ;
        RECT  3.940 0.470 7.165 0.765 ;
        RECT  1.620 3.055 6.520 3.285 ;
        RECT  6.180 2.380 6.520 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.420 3.515 5.760 4.100 ;
        RECT  3.900 3.515 4.240 4.100 ;
        RECT  2.380 3.515 2.720 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  1.065 -0.180 1.405 0.765 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.470 0.685 0.810 ;
        RECT  1.770 1.455 3.960 1.685 ;
        RECT  3.620 1.455 3.960 1.905 ;
        RECT  0.180 0.470 0.410 3.230 ;
        RECT  1.770 1.455 2.000 2.760 ;
        RECT  0.180 2.420 2.000 2.760 ;
        RECT  0.180 2.420 0.520 3.230 ;
    END
END INV_A_NAND4_X4_18_SVT_WB

MACRO INV_A_NAND4_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND4_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.595 1.795 1.030 2.125 ;
        RECT  0.595 1.545 0.935 2.125 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.710 1.770 3.220 2.150 ;
        RECT  2.710 1.520 3.060 2.150 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.620 2.305 2.180 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.260 1.590 1.960 ;
        RECT  1.165 1.260 1.590 1.600 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.977  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.680 2.940 4.200 3.280 ;
        RECT  3.915 0.630 4.200 3.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.960 3.515 4.300 4.100 ;
        RECT  2.440 3.515 2.780 4.100 ;
        RECT  0.920 3.515 1.260 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  0.990 -0.180 1.330 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.360 0.800 3.685 1.030 ;
        RECT  0.360 0.800 0.700 1.290 ;
        RECT  3.450 0.800 3.685 2.710 ;
        RECT  0.360 2.410 3.685 2.710 ;
    END
END INV_A_NAND4_X2_18_SVT_WB

MACRO INV_A_NAND4_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND4_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.210 0.480 1.805 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.225 1.125 2.660 1.590 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.820 2.240 2.250 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.220 1.210 1.790 1.440 ;
        RECT  1.220 1.210 1.560 1.720 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.873  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.520 2.530 3.805 2.870 ;
        RECT  3.575 0.650 3.805 2.870 ;
        RECT  3.350 0.650 3.805 1.030 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.050 3.515 3.675 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.650 3.120 0.880 ;
        RECT  0.180 0.650 0.990 0.980 ;
        RECT  2.890 0.650 3.120 1.730 ;
        RECT  2.890 1.390 3.345 1.730 ;
        RECT  0.710 0.650 0.990 2.720 ;
        RECT  0.180 2.380 0.990 2.720 ;
    END
END INV_A_NAND4_X1_18_SVT_WB

MACRO INV_A_NAND4_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND4_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.760 1.085 2.100 ;
        RECT  0.510 1.370 0.850 2.100 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.260 1.125 2.695 1.590 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.820 2.510 2.135 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.090 1.665 1.590 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.500 2.825 3.790 3.115 ;
        RECT  3.560 0.630 3.790 3.115 ;
        RECT  3.385 0.630 3.790 1.030 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.030 3.515 3.695 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.030 -0.180 1.370 0.400 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.270 0.630 3.155 0.860 ;
        RECT  0.270 0.630 0.610 0.970 ;
        RECT  2.925 0.630 3.155 2.595 ;
        RECT  2.925 2.255 3.330 2.595 ;
        RECT  0.180 2.365 3.330 2.595 ;
        RECT  0.180 2.365 0.520 3.115 ;
    END
END INV_A_NAND4_X0_18_SVT_WB

MACRO INV_A_NAND3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.640 1.640 1.025 2.165 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.980 2.135 4.340 2.365 ;
        RECT  3.930 1.640 4.340 2.365 ;
        RECT  1.980 1.860 2.320 2.365 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.310 2.595 4.940 2.825 ;
        RECT  4.600 1.860 4.940 2.825 ;
        RECT  1.310 1.860 1.650 2.825 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.430  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.020 3.055 5.485 3.395 ;
        RECT  5.170 0.635 5.485 3.395 ;
        RECT  3.020 0.635 5.485 0.865 ;
        RECT  3.020 0.470 3.360 0.865 ;
        RECT  1.500 3.055 5.485 3.285 ;
        RECT  1.500 3.055 1.840 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  2.260 3.515 2.600 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  5.080 -0.180 5.420 0.405 ;
        RECT  1.030 -0.180 1.370 0.880 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.595 0.585 1.410 ;
        RECT  0.180 1.150 3.120 1.410 ;
        RECT  2.780 1.150 3.120 1.905 ;
        RECT  0.180 0.595 0.410 3.215 ;
        RECT  0.180 2.405 0.520 3.215 ;
    END
END INV_A_NAND3_X4_18_SVT_WB

MACRO INV_A_NAND3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.620 2.100 2.235 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.690 1.540 2.150 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.677  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.500 3.045 3.240 3.385 ;
        RECT  3.010 0.550 3.240 3.385 ;
        RECT  2.840 2.410 3.240 3.385 ;
        RECT  2.790 0.550 3.240 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.820 -0.180 1.160 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.040 2.560 1.380 ;
        RECT  2.330 1.840 2.780 2.180 ;
        RECT  2.330 1.040 2.560 2.805 ;
        RECT  0.180 2.465 2.560 2.805 ;
    END
END INV_A_NAND3_X2_18_SVT_WB

MACRO INV_A_NAND3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.815 1.030 2.100 ;
        RECT  0.400 1.600 0.800 2.100 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.610 2.165 2.125 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.165 1.075 1.540 1.620 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.870  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.520 2.880 3.245 3.220 ;
        RECT  3.015 0.510 3.245 3.220 ;
        RECT  2.855 0.510 3.245 0.850 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.725 3.515 1.065 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.940 -0.180 1.280 0.380 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.610 2.625 0.845 ;
        RECT  0.180 0.610 0.520 0.950 ;
        RECT  2.395 0.610 2.625 2.595 ;
        RECT  2.395 2.255 2.785 2.595 ;
        RECT  0.180 2.355 2.785 2.595 ;
        RECT  0.180 2.355 0.520 3.115 ;
    END
END INV_A_NAND3_X1_18_SVT_WB

MACRO INV_A_NAND3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.400 1.815 1.030 2.100 ;
        RECT  0.400 1.600 0.800 2.100 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.610 2.165 2.125 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.165 1.075 1.540 1.620 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.510 2.825 3.245 3.115 ;
        RECT  3.015 0.610 3.245 3.115 ;
        RECT  2.855 0.610 3.245 0.950 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.725 3.515 1.065 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.940 -0.180 1.280 0.380 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.610 2.625 0.845 ;
        RECT  0.180 0.610 0.520 0.950 ;
        RECT  2.395 0.610 2.625 2.595 ;
        RECT  2.395 2.255 2.785 2.595 ;
        RECT  0.180 2.355 2.785 2.595 ;
        RECT  0.180 2.355 0.520 3.115 ;
    END
END INV_A_NAND3_X0_18_SVT_WB

MACRO INV_A_NAND2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.160 0.600 1.960 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.840 2.135 6.630 2.365 ;
        RECT  6.220 1.800 6.630 2.365 ;
        RECT  3.980 1.915 4.320 2.365 ;
        RECT  1.840 1.915 2.180 2.365 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.618  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 2.595 7.165 2.935 ;
        RECT  6.860 0.995 7.165 2.935 ;
        RECT  2.780 0.995 7.165 1.225 ;
        RECT  6.115 2.595 6.505 3.425 ;
        RECT  5.420 0.470 5.760 1.225 ;
        RECT  4.820 2.595 5.160 3.350 ;
        RECT  3.500 2.595 3.840 3.405 ;
        RECT  2.060 2.595 7.165 2.835 ;
        RECT  2.780 0.515 3.120 1.225 ;
        RECT  2.060 2.595 2.400 3.405 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  2.780 3.065 3.120 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.760 -0.180 7.100 0.765 ;
        RECT  4.220 -0.180 4.560 0.765 ;
        RECT  1.630 -0.180 1.970 0.810 ;
        RECT  0.190 -0.180 0.530 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.910 1.455 5.540 1.685 ;
        RECT  2.540 1.455 2.880 1.905 ;
        RECT  5.200 1.455 5.540 1.905 ;
        RECT  0.910 0.470 1.250 3.190 ;
        RECT  0.740 2.380 1.250 3.190 ;
    END
END INV_A_NAND2_X8_18_SVT_WB

MACRO INV_A_NAND2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.336  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.680 0.570 2.150 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.550 1.820 3.345 2.200 ;
        RECT  1.260 2.135 2.890 2.365 ;
        RECT  1.260 1.860 1.600 2.365 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.809  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.500 2.595 3.805 2.935 ;
        RECT  3.575 0.645 3.805 2.935 ;
        RECT  2.150 0.645 3.805 0.875 ;
        RECT  2.820 2.595 3.220 3.405 ;
        RECT  2.150 0.470 2.490 0.875 ;
        RECT  1.500 2.595 1.840 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.340 -0.180 3.680 0.415 ;
        RECT  0.940 -0.180 1.280 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.535 0.520 1.440 ;
        RECT  0.180 1.105 2.320 1.440 ;
        RECT  0.800 1.105 2.320 1.445 ;
        RECT  1.980 1.105 2.320 1.905 ;
        RECT  0.800 1.105 1.030 2.720 ;
        RECT  0.180 2.380 1.030 2.720 ;
    END
END INV_A_NAND2_X4_18_SVT_WB

MACRO INV_A_NAND2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.210 1.160 1.590 ;
        RECT  0.425 1.620 0.930 1.960 ;
        RECT  0.700 1.210 0.930 1.960 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.160 1.820 1.590 2.290 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.356  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.505 3.045 2.660 3.285 ;
        RECT  2.290 0.470 2.660 3.285 ;
        RECT  1.505 3.045 1.845 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.265 3.515 2.605 4.100 ;
        RECT  0.745 3.515 1.085 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.350 -0.180 1.165 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.185 0.750 2.060 0.980 ;
        RECT  0.185 0.750 0.470 1.335 ;
        RECT  0.185 2.410 0.525 2.750 ;
        RECT  1.820 0.750 2.060 2.750 ;
        RECT  0.185 2.520 2.060 2.750 ;
    END
END INV_A_NAND2_X2_18_SVT_WB

MACRO INV_A_NAND2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.450 1.725 0.980 2.205 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.105 1.605 1.570 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.562  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.520 2.930 2.660 3.270 ;
        RECT  2.295 0.540 2.660 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.280 3.500 2.620 4.100 ;
        RECT  0.760 3.515 1.100 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.050 -0.180 1.390 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.645 2.065 0.875 ;
        RECT  0.180 0.645 0.520 0.985 ;
        RECT  1.740 2.255 2.065 2.700 ;
        RECT  1.835 0.645 2.065 2.700 ;
        RECT  0.200 2.470 2.065 2.700 ;
        RECT  0.200 2.470 0.540 3.115 ;
    END
END INV_A_NAND2_X1_18_SVT_WB

MACRO INV_A_NAND2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.620 0.670 2.350 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.830 1.745 9.965 2.200 ;
        RECT  2.000 2.180 9.170 2.410 ;
        RECT  7.020 1.915 7.360 2.410 ;
        RECT  4.620 1.915 4.960 2.410 ;
        RECT  2.000 1.915 2.340 2.410 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.427  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.640 10.500 2.870 ;
        RECT  10.195 1.050 10.500 2.870 ;
        RECT  8.680 1.050 10.500 1.420 ;
        RECT  9.400 2.640 9.740 3.455 ;
        RECT  7.980 2.640 9.740 2.980 ;
        RECT  2.940 0.985 9.020 1.225 ;
        RECT  8.680 0.610 9.020 1.420 ;
        RECT  7.980 2.640 8.320 3.450 ;
        RECT  2.220 2.640 9.740 2.880 ;
        RECT  6.540 2.640 6.880 3.450 ;
        RECT  5.100 2.640 5.440 3.450 ;
        RECT  3.660 2.640 4.000 3.450 ;
        RECT  2.220 2.640 4.000 2.980 ;
        RECT  2.940 0.470 3.290 1.225 ;
        RECT  2.220 2.640 2.560 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  10.120 3.100 10.460 4.100 ;
        RECT  7.260 3.110 7.600 4.100 ;
        RECT  5.820 3.110 6.160 4.100 ;
        RECT  4.380 3.110 4.720 4.100 ;
        RECT  0.185 2.630 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  10.120 -0.180 10.460 0.810 ;
        RECT  7.260 -0.180 7.600 0.755 ;
        RECT  4.380 -0.180 4.720 0.755 ;
        RECT  1.620 -0.180 1.960 0.810 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 1.455 8.270 1.685 ;
        RECT  2.700 1.455 3.040 1.950 ;
        RECT  5.600 1.455 5.940 1.950 ;
        RECT  8.045 1.620 8.550 1.950 ;
        RECT  0.900 0.470 1.240 3.450 ;
    END
END INV_A_NAND2_X12_18_SVT_WB

MACRO INV_A_NAND2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_NAND2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN AN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.445 1.710 0.980 2.190 ;
        END
    END AN
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.105 1.605 1.550 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.670 2.465 2.660 2.695 ;
        RECT  2.295 0.645 2.660 2.695 ;
        RECT  1.520 2.995 1.900 3.280 ;
        RECT  1.670 2.465 1.900 3.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  2.280 2.925 2.620 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.050 -0.180 1.390 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.645 2.065 0.875 ;
        RECT  0.180 0.645 0.520 0.985 ;
        RECT  1.835 0.645 2.065 2.235 ;
        RECT  1.210 1.850 2.065 2.235 ;
        RECT  1.210 1.850 1.440 2.760 ;
        RECT  0.180 2.420 1.440 2.760 ;
        RECT  0.180 2.420 0.520 3.280 ;
    END
END INV_A_NAND2_X0_18_SVT_WB

MACRO INV_A_INV_B_OAI22_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_INV_B_OAI22_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.875 1.725 4.455 2.150 ;
        RECT  3.875 1.260 4.215 2.150 ;
        RECT  3.675 1.260 4.215 1.600 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.725 1.655 6.300 2.215 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.675 0.760 2.190 ;
        END
    END B0
    PIN B1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.670 2.325 2.185 ;
        END
    END B1N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.468  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.115 2.950 8.265 3.285 ;
        RECT  7.900 1.085 8.265 3.285 ;
        RECT  5.775 1.085 8.265 1.425 ;
        RECT  2.115 2.420 2.455 3.285 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.630 3.515 7.970 4.100 ;
        RECT  4.960 3.515 5.300 4.100 ;
        RECT  3.340 3.515 3.680 4.100 ;
        RECT  0.920 3.110 1.260 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  3.630 -0.180 3.970 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 0.505 0.540 1.315 ;
        RECT  0.200 1.085 3.445 1.315 ;
        RECT  3.105 1.085 3.445 1.960 ;
        RECT  1.160 1.085 1.500 2.760 ;
        RECT  0.200 2.420 1.500 2.760 ;
        RECT  0.200 2.420 0.540 3.230 ;
        RECT  4.445 1.100 5.470 1.440 ;
        RECT  6.575 1.655 7.670 2.025 ;
        RECT  5.170 1.100 5.470 2.720 ;
        RECT  4.100 2.380 5.470 2.720 ;
        RECT  6.575 1.655 6.915 2.720 ;
        RECT  4.100 2.480 6.915 2.720 ;
        RECT  5.000 0.470 5.340 0.855 ;
        RECT  7.880 0.515 8.220 0.855 ;
        RECT  1.550 0.580 8.220 0.855 ;
    END
END INV_A_INV_B_OAI22_X4_18_SVT_WB

MACRO INV_A_INV_B_OAI22_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_INV_B_OAI22_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.060 0.505 2.725 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.615 4.390 2.150 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.715 1.740 2.100 ;
        END
    END B0
    PIN B1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.435 1.210 3.780 1.980 ;
        END
    END B1N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.620 1.105 4.975 1.440 ;
        RECT  3.915 2.380 4.850 2.720 ;
        RECT  4.620 1.105 4.850 2.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.540 2.380 5.825 4.100 ;
        RECT  1.255 3.525 2.825 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  3.155 -0.180 3.495 0.405 ;
        RECT  0.975 -0.180 1.315 0.825 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.695 0.555 2.030 1.365 ;
        RECT  1.970 1.135 2.200 2.720 ;
        RECT  1.970 1.860 3.090 2.200 ;
        RECT  1.970 1.860 2.310 2.720 ;
        RECT  0.265 0.645 0.595 1.740 ;
        RECT  0.265 1.510 0.980 1.740 ;
        RECT  5.080 1.825 5.455 2.165 ;
        RECT  0.735 1.510 0.980 3.295 ;
        RECT  5.080 1.825 5.310 3.295 ;
        RECT  0.255 2.955 5.310 3.295 ;
        RECT  2.395 0.535 2.735 0.875 ;
        RECT  3.915 0.535 5.695 0.875 ;
        RECT  2.395 0.635 5.695 0.875 ;
        RECT  5.355 0.535 5.695 1.440 ;
    END
END INV_A_INV_B_OAI22_X2_18_SVT_WB

MACRO INV_A_INV_B_OAI22_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_INV_B_OAI22_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.050 0.980 1.960 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.820 4.695 2.150 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.385 1.670 2.150 2.100 ;
        END
    END B0
    PIN B1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.120 3.950 1.590 ;
        END
    END B1N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.631  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.130 2.380 5.250 2.820 ;
        RECT  4.925 1.100 5.250 2.820 ;
        RECT  4.850 1.100 5.250 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.570 2.535 5.950 4.100 ;
        RECT  2.980 2.535 3.320 4.100 ;
        RECT  0.905 2.910 1.245 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  3.330 -0.180 3.670 0.350 ;
        RECT  0.970 -0.180 1.325 0.820 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.185 0.640 0.470 3.250 ;
        RECT  0.185 2.340 2.195 2.680 ;
        RECT  0.185 2.340 0.525 3.250 ;
        RECT  1.795 0.615 2.135 1.440 ;
        RECT  1.795 1.100 2.735 1.440 ;
        RECT  2.435 1.100 2.735 3.250 ;
        RECT  1.625 2.910 2.735 3.250 ;
        RECT  2.570 0.580 5.970 0.870 ;
        RECT  5.570 0.580 5.970 1.335 ;
    END
END INV_A_INV_B_OAI22_X1_18_SVT_WB

MACRO INV_A_INV_B_OAI22_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_INV_B_OAI22_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.260 1.030 1.600 ;
        RECT  0.650 1.260 0.940 1.930 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.555 4.405 2.150 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.170 1.790 1.665 2.130 ;
        RECT  1.380 1.275 1.665 2.130 ;
        END
    END B0
    PIN B1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.495 3.830 2.100 ;
        END
    END B1N
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.930 2.540 4.865 2.880 ;
        RECT  4.635 0.925 4.865 2.880 ;
        RECT  4.360 0.925 4.865 1.265 ;
        RECT  3.930 2.380 4.390 2.880 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  5.095 2.395 5.420 4.100 ;
        RECT  2.815 2.395 3.120 4.100 ;
        RECT  0.900 2.940 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  2.790 -0.180 3.130 0.405 ;
        RECT  0.900 -0.180 1.240 1.030 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.705 0.520 1.045 ;
        RECT  0.180 0.705 0.420 3.280 ;
        RECT  0.180 2.365 2.125 2.705 ;
        RECT  0.180 2.365 0.520 3.280 ;
        RECT  1.620 0.705 2.125 1.045 ;
        RECT  1.895 0.705 2.125 2.135 ;
        RECT  1.895 1.795 2.900 2.135 ;
        RECT  2.355 1.795 2.585 3.280 ;
        RECT  1.620 2.940 2.585 3.280 ;
        RECT  3.640 0.410 5.420 0.695 ;
        RECT  3.640 0.410 3.980 1.265 ;
        RECT  2.355 0.925 3.980 1.265 ;
        RECT  5.095 0.410 5.420 1.265 ;
    END
END INV_A_INV_B_OAI22_X0_18_SVT_WB

MACRO INV_A_AOI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AOI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.210 2.700 1.960 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.100 0.500 1.665 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.620 1.670 2.155 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.305 2.545 7.645 3.385 ;
        RECT  5.985 1.055 7.645 1.350 ;
        RECT  7.305 0.535 7.645 1.350 ;
        RECT  5.985 2.545 7.645 2.940 ;
        RECT  6.780 1.055 7.155 2.940 ;
        RECT  5.985 0.590 6.335 1.350 ;
        RECT  5.985 2.545 6.325 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  5.220 3.570 5.560 4.100 ;
        RECT  1.105 3.515 1.445 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  5.220 -0.180 5.560 0.350 ;
        RECT  3.625 -0.180 4.010 1.390 ;
        RECT  1.105 -0.180 1.445 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.345 0.535 0.685 0.870 ;
        RECT  0.345 0.640 3.160 0.870 ;
        RECT  2.930 0.640 3.160 1.960 ;
        RECT  2.930 1.620 3.405 1.960 ;
        RECT  0.730 0.640 0.960 2.720 ;
        RECT  0.340 2.380 0.960 2.720 ;
        RECT  1.865 3.045 3.645 3.385 ;
        RECT  4.050 1.750 4.780 2.085 ;
        RECT  1.900 1.100 2.150 2.720 ;
        RECT  4.050 1.750 4.385 2.720 ;
        RECT  1.900 2.380 4.385 2.720 ;
        RECT  4.660 0.905 5.345 1.160 ;
        RECT  5.010 0.905 5.345 2.670 ;
        RECT  5.010 1.620 6.525 1.960 ;
        RECT  5.010 1.620 5.350 2.670 ;
        RECT  4.660 2.405 5.350 2.670 ;
    END
END INV_A_AOI21_X8_18_SVT_WB

MACRO INV_A_AOI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AOI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.205 1.510 2.730 2.130 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.196  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.630 0.480 2.205 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.535 2.910 1.430 3.220 ;
        RECT  1.170 1.620 1.430 3.220 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.080 2.565 6.020 2.895 ;
        RECT  5.720 1.015 6.020 2.895 ;
        RECT  5.080 1.015 6.020 1.365 ;
        RECT  5.080 2.565 5.435 3.385 ;
        RECT  5.080 0.535 5.405 1.365 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.320 3.515 4.660 4.100 ;
        RECT  0.860 3.515 1.200 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.320 -0.180 4.660 0.405 ;
        RECT  3.115 -0.180 3.400 0.820 ;
        RECT  0.860 -0.180 1.200 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.685 0.640 2.885 0.870 ;
        RECT  2.655 0.640 2.885 1.280 ;
        RECT  2.655 1.050 3.285 1.280 ;
        RECT  0.685 0.640 0.940 1.365 ;
        RECT  0.180 1.010 0.940 1.365 ;
        RECT  2.960 1.050 3.285 1.960 ;
        RECT  0.710 0.640 0.940 2.665 ;
        RECT  0.175 2.435 0.940 2.665 ;
        RECT  1.675 3.045 3.400 3.385 ;
        RECT  1.655 1.100 1.975 1.455 ;
        RECT  3.710 1.800 4.305 2.180 ;
        RECT  1.745 1.100 1.975 2.665 ;
        RECT  2.375 2.360 3.940 2.590 ;
        RECT  3.710 1.800 3.940 2.590 ;
        RECT  1.745 2.435 2.690 2.665 ;
        RECT  3.760 1.095 4.100 1.485 ;
        RECT  3.760 1.255 4.850 1.485 ;
        RECT  4.535 1.625 5.245 1.965 ;
        RECT  4.535 1.255 4.850 3.105 ;
        RECT  3.760 2.820 4.850 3.105 ;
    END
END INV_A_AOI21_X4_18_SVT_WB

MACRO INV_A_AOI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AOI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.210 2.700 1.960 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.100 0.500 1.665 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.620 1.670 2.155 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.900 2.380 3.305 2.720 ;
        RECT  1.900 1.100 2.150 2.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.105 3.515 1.445 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.390 -0.180 3.675 1.390 ;
        RECT  1.105 -0.180 1.445 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.345 0.535 0.685 0.870 ;
        RECT  0.345 0.640 3.160 0.870 ;
        RECT  2.930 0.640 3.160 1.960 ;
        RECT  2.930 1.620 3.405 1.960 ;
        RECT  0.730 0.640 0.960 2.720 ;
        RECT  0.340 2.380 0.960 2.720 ;
        RECT  1.865 3.045 3.645 3.385 ;
    END
END INV_A_AOI21_X2_18_SVT_WB

MACRO INV_A_AOI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AOI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.460 2.130 2.170 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.595 0.980 2.150 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.175 1.580 2.690 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.360 0.635 2.770 0.985 ;
        RECT  2.200 2.400 2.590 2.740 ;
        RECT  2.360 0.635 2.590 2.740 ;
        RECT  1.720 0.635 2.770 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.840 3.515 1.180 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.000 -0.180 1.340 0.945 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.635 0.620 0.975 ;
        RECT  0.115 0.635 0.345 3.200 ;
        RECT  0.115 2.555 0.620 3.200 ;
        RECT  2.820 1.880 3.160 3.200 ;
        RECT  0.115 2.970 3.160 3.200 ;
    END
END INV_A_AOI21_X1_18_SVT_WB

MACRO INV_A_AOI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AOI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.795 1.540 2.200 2.160 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.820 1.070 2.100 ;
        RECT  0.575 1.430 0.860 2.100 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.185 1.070 1.565 1.605 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.200 2.390 2.660 2.720 ;
        RECT  2.430 0.535 2.660 2.720 ;
        RECT  2.380 0.535 2.660 1.185 ;
        RECT  1.720 0.535 2.660 0.875 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.840 3.515 1.180 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.000 -0.180 1.340 0.840 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.535 0.620 0.875 ;
        RECT  0.115 0.535 0.345 3.180 ;
        RECT  0.115 2.775 0.620 3.180 ;
        RECT  2.890 1.860 3.195 3.180 ;
        RECT  0.115 2.950 3.195 3.180 ;
    END
END INV_A_AOI21_X0_18_SVT_WB

MACRO INV_A_AO22_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AO22_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.840 2.100 2.780 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.950 1.715 4.385 2.180 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 0.650 1.375 1.960 ;
        RECT  0.700 0.650 1.375 1.100 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.180 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.080 2.380 5.460 3.300 ;
        RECT  5.135 0.470 5.460 3.300 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  3.850 3.515 4.660 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  2.760 -0.180 3.100 0.400 ;
        RECT  0.180 -0.180 0.470 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.415 0.520 3.350 ;
        RECT  0.180 3.010 3.350 3.350 ;
        RECT  3.470 1.100 3.810 1.440 ;
        RECT  3.470 1.100 3.720 2.200 ;
        RECT  3.000 1.860 3.720 2.200 ;
        RECT  3.490 1.100 3.720 2.750 ;
        RECT  3.490 2.410 4.050 2.750 ;
        RECT  1.605 0.630 4.905 0.870 ;
        RECT  1.605 0.630 2.630 0.970 ;
        RECT  1.605 0.630 1.910 1.440 ;
        RECT  4.620 0.630 4.905 1.960 ;
        RECT  2.330 0.630 2.630 2.720 ;
    END
END INV_A_AO22_X4_18_SVT_WB

MACRO INV_A_AO22_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AO22_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.860 2.150 2.710 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.000 1.040 4.340 1.740 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.095 1.640 1.640 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.520 0.980 2.150 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.080 2.420 5.460 3.385 ;
        RECT  5.230 0.570 5.460 3.385 ;
        RECT  5.080 0.570 5.460 1.455 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.320 3.515 4.660 4.100 ;
        RECT  0.860 3.515 1.200 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.360 -0.180 4.700 0.810 ;
        RECT  2.920 -0.180 3.260 0.915 ;
        RECT  0.300 -0.180 0.640 0.915 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.300 2.775 0.640 3.195 ;
        RECT  0.300 2.965 1.960 3.195 ;
        RECT  1.620 2.965 1.960 3.345 ;
        RECT  3.540 0.470 3.980 0.810 ;
        RECT  3.170 1.210 3.770 1.550 ;
        RECT  3.540 0.470 3.770 2.720 ;
        RECT  3.540 2.380 4.100 2.720 ;
        RECT  1.800 0.575 2.690 0.925 ;
        RECT  4.620 1.860 5.000 2.200 ;
        RECT  2.380 0.575 2.690 3.285 ;
        RECT  4.620 1.860 4.850 3.285 ;
        RECT  2.380 2.950 4.850 3.285 ;
    END
END INV_A_AO22_X2_18_SVT_WB

MACRO INV_A_AO22_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AO22_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.140 2.245 1.620 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.780 4.260 2.170 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.260 1.590 2.120 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.185 0.980 1.900 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.105 0.595 5.460 2.765 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.320 3.515 4.660 4.100 ;
        RECT  0.940 3.005 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  2.975 -0.180 3.300 0.880 ;
        RECT  0.180 -0.180 0.520 0.910 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.535 2.040 2.775 ;
        RECT  0.180 2.535 0.520 2.875 ;
        RECT  1.700 2.535 2.040 2.875 ;
        RECT  3.680 0.690 4.020 1.495 ;
        RECT  2.955 1.165 4.020 1.495 ;
        RECT  2.955 1.165 3.220 2.720 ;
        RECT  2.955 2.400 4.020 2.720 ;
        RECT  1.700 0.570 2.725 0.910 ;
        RECT  2.475 0.570 2.725 3.180 ;
        RECT  4.590 1.715 4.875 3.180 ;
        RECT  2.475 2.950 4.875 3.180 ;
    END
END INV_A_AO22_X1_18_SVT_WB

MACRO INV_A_AO22_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN INV_A_AO22_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.140 2.245 1.620 ;
        END
    END A0
    PIN A1N
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.805 4.260 2.190 ;
        END
    END A1N
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.260 1.590 2.120 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.620 1.185 0.980 1.900 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.105 0.680 5.460 2.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.320 3.515 4.660 4.100 ;
        RECT  0.940 3.005 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  2.955 -0.180 3.300 0.875 ;
        RECT  0.180 -0.180 0.520 0.910 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.535 2.040 2.775 ;
        RECT  0.180 2.535 0.520 2.875 ;
        RECT  1.700 2.535 2.040 2.875 ;
        RECT  3.680 0.690 4.020 1.490 ;
        RECT  2.955 1.165 4.020 1.490 ;
        RECT  2.955 1.165 3.220 2.720 ;
        RECT  2.955 2.430 4.020 2.720 ;
        RECT  1.700 0.570 2.725 0.910 ;
        RECT  2.475 0.570 2.725 3.180 ;
        RECT  4.590 1.715 4.875 3.180 ;
        RECT  2.475 2.950 4.875 3.180 ;
    END
END INV_A_AO22_X0_18_SVT_WB

MACRO INVP2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.003  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.510 3.790 2.100 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.221  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.755 2.330 4.250 2.720 ;
        RECT  4.020 0.535 4.250 2.720 ;
        RECT  0.755 1.050 4.250 1.280 ;
        RECT  3.825 0.535 4.250 1.280 ;
        RECT  2.275 0.535 2.660 1.280 ;
        RECT  2.075 2.330 2.445 3.085 ;
        RECT  0.755 0.750 1.095 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.960 3.515 4.300 4.100 ;
        RECT  0.180 3.515 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.035 -0.180 3.375 0.820 ;
        RECT  1.515 -0.180 1.855 0.820 ;
        END
    END VSS
END INVP2_X8_18_SVT_WB

MACRO INVP2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.672  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.565 3.155 1.905 ;
        RECT  0.575 1.565 1.030 2.100 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.112  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.080 2.555 3.740 3.310 ;
        RECT  3.400 0.590 3.740 3.310 ;
        RECT  0.330 1.105 3.740 1.335 ;
        RECT  2.080 2.140 2.420 3.310 ;
        RECT  0.330 1.100 2.200 1.335 ;
        RECT  1.860 0.805 2.200 1.335 ;
        RECT  0.760 2.555 3.740 2.895 ;
        RECT  0.330 0.805 0.670 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.180 3.515 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  2.640 -0.180 2.980 0.875 ;
        RECT  1.100 -0.180 1.440 0.870 ;
        END
    END VSS
END INVP2_X6_18_SVT_WB

MACRO INVP2_X5_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.225 1.620 1.395 2.100 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.611  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.870 3.780 3.450 ;
        RECT  0.760 2.640 3.780 2.980 ;
        RECT  3.400 0.870 3.780 2.980 ;
        RECT  2.080 2.640 2.420 3.395 ;
        RECT  2.005 1.100 2.300 2.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.180 3.515 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  2.680 -0.180 3.020 1.220 ;
        RECT  1.240 -0.180 1.580 1.240 ;
        END
    END VSS
END INVP2_X5_18_SVT_WB

MACRO INVP2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.206  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.235 1.620 1.875 2.365 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.809  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.640 2.525 3.450 ;
        RECT  2.105 0.575 2.525 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 2.695 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.780 -0.180 3.120 1.330 ;
        RECT  1.340 -0.180 1.680 1.385 ;
        END
    END VSS
END INVP2_X4_18_SVT_WB

MACRO INVP2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.904  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 1.495 1.415 2.200 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.597  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 2.695 2.620 3.450 ;
        RECT  0.900 2.695 2.620 3.220 ;
        RECT  1.735 0.975 2.015 3.220 ;
        RECT  1.615 0.975 2.015 1.315 ;
        RECT  0.900 2.695 1.240 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.695 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.280 -0.180 2.620 1.045 ;
        RECT  0.840 -0.180 1.180 1.265 ;
        END
    END VSS
END INVP2_X3_18_SVT_WB

MACRO INVP2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.603  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.205 1.780 1.905 2.120 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.125  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 2.435 1.240 3.270 ;
        RECT  0.700 1.815 0.930 3.270 ;
        RECT  0.430 0.685 0.770 2.065 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.620 2.435 1.960 4.100 ;
        RECT  0.180 2.380 0.470 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.160 -0.180 1.480 1.440 ;
        END
    END VSS
END INVP2_X2_18_SVT_WB

MACRO INVP2_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 7.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.715 1.245 8.950 1.585 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 11.607  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.360 2.630 14.700 3.385 ;
        RECT  9.505 0.680 14.700 1.020 ;
        RECT  11.220 2.630 14.700 2.970 ;
        RECT  12.740 2.630 13.080 3.330 ;
        RECT  11.220 2.630 11.560 3.330 ;
        RECT  8.260 2.630 14.700 2.895 ;
        RECT  9.505 0.680 10.400 2.895 ;
        RECT  9.780 0.680 10.120 3.330 ;
        RECT  8.260 2.630 10.120 2.970 ;
        RECT  0.900 0.680 14.700 1.015 ;
        RECT  8.260 2.630 8.600 3.395 ;
        RECT  0.900 2.630 14.700 2.880 ;
        RECT  6.820 2.630 7.160 3.330 ;
        RECT  5.300 2.630 7.160 2.970 ;
        RECT  5.300 2.630 5.640 3.330 ;
        RECT  3.860 2.630 4.200 3.330 ;
        RECT  2.340 2.630 4.200 2.970 ;
        RECT  2.340 2.630 2.680 3.330 ;
        RECT  0.900 2.630 4.200 2.945 ;
        RECT  0.900 2.630 1.240 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.120 4.100 ;
        RECT  13.500 3.320 13.840 4.100 ;
        RECT  11.980 3.515 12.320 4.100 ;
        RECT  10.500 3.125 10.840 4.100 ;
        RECT  9.020 3.515 9.360 4.100 ;
        RECT  7.540 3.110 7.880 4.100 ;
        RECT  6.060 3.515 6.400 4.100 ;
        RECT  4.580 3.110 4.920 4.100 ;
        RECT  3.100 3.515 3.440 4.100 ;
        RECT  1.620 3.175 1.960 4.100 ;
        RECT  0.180 2.685 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.120 0.180 ;
        RECT  12.160 -0.180 12.500 0.405 ;
        RECT  9.200 -0.180 9.540 0.410 ;
        RECT  6.240 -0.180 6.580 0.405 ;
        RECT  3.280 -0.180 3.620 0.410 ;
        RECT  0.180 -0.180 0.520 1.065 ;
        END
    END VSS
END INVP2_X24_18_SVT_WB

MACRO INVP2_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.805  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.685 1.245 6.365 1.585 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.109  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.240 2.575 11.580 3.385 ;
        RECT  0.920 0.685 11.580 1.015 ;
        RECT  0.920 2.575 11.580 2.880 ;
        RECT  9.800 2.575 10.140 3.385 ;
        RECT  8.280 2.575 10.140 2.915 ;
        RECT  8.280 2.575 8.620 3.385 ;
        RECT  6.840 0.685 7.595 2.880 ;
        RECT  6.840 0.685 7.180 3.385 ;
        RECT  2.360 2.575 7.180 2.915 ;
        RECT  5.320 2.575 5.660 3.385 ;
        RECT  3.880 2.575 4.220 3.385 ;
        RECT  2.360 2.575 2.700 3.385 ;
        RECT  0.920 2.420 1.260 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  10.520 3.110 10.860 4.100 ;
        RECT  9.040 3.515 9.380 4.100 ;
        RECT  7.560 3.110 7.900 4.100 ;
        RECT  6.080 3.515 6.420 4.100 ;
        RECT  4.600 3.145 4.940 4.100 ;
        RECT  3.120 3.515 3.460 4.100 ;
        RECT  1.640 3.110 1.980 4.100 ;
        RECT  0.200 2.420 0.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  9.040 -0.180 9.380 0.350 ;
        RECT  6.080 -0.180 6.420 0.410 ;
        RECT  3.120 -0.180 3.460 0.410 ;
        RECT  0.200 -0.180 0.540 1.065 ;
        END
    END VSS
END INVP2_X20_18_SVT_WB

MACRO INVP2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.301  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.165 0.920 1.590 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.804  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 0.645 1.540 3.175 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  0.430 2.640 0.770 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  0.430 -0.180 0.770 0.880 ;
        END
    END VSS
END INVP2_X1_18_SVT_WB

MACRO INVP2_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.430 1.490 4.560 2.100 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.705  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.880 2.640 8.220 3.450 ;
        RECT  0.900 0.995 8.220 1.225 ;
        RECT  7.880 0.730 8.220 1.225 ;
        RECT  0.900 2.640 8.220 2.880 ;
        RECT  6.440 2.640 6.780 3.450 ;
        RECT  5.120 0.700 6.780 1.225 ;
        RECT  5.120 2.640 6.780 2.980 ;
        RECT  4.835 0.995 5.720 2.880 ;
        RECT  5.120 0.700 5.460 3.450 ;
        RECT  3.680 2.640 4.020 3.450 ;
        RECT  2.340 0.730 4.020 1.225 ;
        RECT  2.340 2.640 4.020 2.980 ;
        RECT  2.340 2.640 2.680 3.450 ;
        RECT  0.900 2.640 1.240 3.450 ;
        RECT  0.900 0.730 1.240 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.160 3.110 7.500 4.100 ;
        RECT  4.400 3.110 4.740 4.100 ;
        RECT  1.620 3.110 1.960 4.100 ;
        RECT  0.180 2.420 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.160 -0.180 7.500 0.765 ;
        RECT  4.400 -0.180 4.740 0.765 ;
        RECT  1.620 -0.180 1.960 0.765 ;
        RECT  0.180 -0.180 0.520 1.070 ;
        END
    END VSS
END INVP2_X16_18_SVT_WB

MACRO INVP2_X14_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X14_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.595  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.085 1.260 3.665 1.660 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.631  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.895 0.985 7.070 1.215 ;
        RECT  6.730 0.690 7.070 1.215 ;
        RECT  6.190 2.225 6.530 2.930 ;
        RECT  0.900 2.225 6.530 2.455 ;
        RECT  0.900 0.970 5.630 1.030 ;
        RECT  5.290 0.470 5.630 1.215 ;
        RECT  4.860 2.225 5.200 3.395 ;
        RECT  3.895 0.970 4.440 2.455 ;
        RECT  0.900 0.690 4.190 1.030 ;
        RECT  3.540 2.225 3.880 2.930 ;
        RECT  2.210 2.225 2.560 3.395 ;
        RECT  0.900 2.225 1.240 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.760 3.515 7.100 4.100 ;
        RECT  2.980 3.515 3.320 4.100 ;
        RECT  0.180 2.695 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.010 -0.180 6.350 0.755 ;
        RECT  4.570 -0.180 4.910 0.740 ;
        RECT  3.090 -0.180 3.430 0.460 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
END INVP2_X14_18_SVT_WB

MACRO INVP2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.179  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 1.510 3.350 2.100 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.972  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.880 2.770 6.540 3.110 ;
        RECT  5.380 0.740 5.720 1.265 ;
        RECT  3.940 1.035 5.720 1.265 ;
        RECT  4.880 2.105 5.220 3.385 ;
        RECT  3.580 2.370 5.220 2.915 ;
        RECT  3.580 1.050 4.340 2.915 ;
        RECT  3.940 0.535 4.280 2.915 ;
        RECT  0.900 2.575 5.220 2.915 ;
        RECT  0.900 1.050 4.340 1.280 ;
        RECT  2.420 0.740 2.760 1.280 ;
        RECT  2.240 2.575 2.580 3.385 ;
        RECT  0.900 2.380 1.240 3.190 ;
        RECT  0.900 0.740 1.240 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  5.640 3.515 6.450 4.100 ;
        RECT  3.000 3.515 3.340 4.100 ;
        RECT  0.180 2.380 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  6.100 -0.180 6.440 0.930 ;
        RECT  4.660 -0.180 5.000 0.805 ;
        RECT  3.180 -0.180 3.520 0.820 ;
        RECT  1.660 -0.180 2.000 0.820 ;
        RECT  0.180 -0.180 0.520 0.860 ;
        END
    END VSS
END INVP2_X12_18_SVT_WB

MACRO INVP2_X10_18_SVT_WB
    CLASS CORE ;
    FOREIGN INVP2_X10_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.857  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.595 1.510 4.275 2.105 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.600  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.520 2.640 5.180 3.395 ;
        RECT  4.860 0.535 5.180 3.395 ;
        RECT  4.840 1.050 5.180 3.395 ;
        RECT  0.300 1.050 5.180 1.280 ;
        RECT  3.340 0.535 3.800 1.280 ;
        RECT  0.760 2.640 5.180 2.895 ;
        RECT  2.080 2.640 2.420 3.395 ;
        RECT  1.820 0.755 2.160 1.280 ;
        RECT  0.760 2.640 2.420 2.980 ;
        RECT  0.300 0.760 0.640 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.640 2.575 5.980 4.100 ;
        RECT  2.800 3.125 3.140 4.100 ;
        RECT  0.180 3.515 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  5.600 -0.180 5.940 0.820 ;
        RECT  4.100 -0.180 4.440 0.820 ;
        RECT  2.580 -0.180 2.920 0.820 ;
        RECT  1.060 -0.180 1.400 0.820 ;
        END
    END VSS
END INVP2_X10_18_SVT_WB

MACRO HOLD_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN HOLD_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Q
        DIRECTION INOUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.105 1.625 2.200 ;
        RECT  0.190 1.105 1.625 1.410 ;
        RECT  0.190 0.470 0.530 1.410 ;
        RECT  0.190 0.470 0.495 2.755 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.950 2.900 1.290 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.950 -0.180 1.290 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.710 0.535 2.110 0.875 ;
        RECT  0.725 1.640 1.010 2.670 ;
        RECT  0.725 2.430 2.110 2.670 ;
        RECT  1.855 0.535 2.110 3.385 ;
        RECT  1.710 2.430 2.110 3.385 ;
    END
END HOLD_X1_18_SVT_WB

MACRO HA1_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN HA1_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.355 2.135 6.450 2.365 ;
        RECT  6.110 1.860 6.450 2.365 ;
        RECT  3.355 1.770 3.780 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.050 1.620 5.060 1.905 ;
        RECT  4.050 1.210 4.590 1.905 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.420 2.665 3.230 ;
        RECT  2.175 0.580 2.665 1.390 ;
        RECT  2.175 0.580 2.405 2.760 ;
        RECT  0.900 1.760 2.405 2.100 ;
        RECT  0.900 0.635 1.240 3.175 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.360 0.550 9.700 3.190 ;
        RECT  7.965 1.985 9.700 2.325 ;
        RECT  7.965 0.535 8.260 3.245 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  10.120 2.490 10.460 4.100 ;
        RECT  8.640 2.710 8.980 4.100 ;
        RECT  7.160 3.515 7.500 4.100 ;
        RECT  4.500 3.110 5.540 4.100 ;
        RECT  3.060 3.110 3.400 4.100 ;
        RECT  1.620 2.640 1.945 4.100 ;
        RECT  0.180 2.695 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  10.080 -0.180 10.420 1.250 ;
        RECT  8.640 -0.180 8.980 1.290 ;
        RECT  7.160 -0.180 7.500 0.820 ;
        RECT  3.060 -0.180 3.360 0.810 ;
        RECT  1.620 -0.180 1.945 1.390 ;
        RECT  0.180 -0.180 0.520 1.335 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  4.910 0.530 6.690 0.875 ;
        RECT  4.910 0.530 5.250 1.230 ;
        RECT  3.590 0.695 4.550 0.980 ;
        RECT  3.590 0.695 3.820 1.540 ;
        RECT  2.895 1.200 3.820 1.540 ;
        RECT  2.635 1.620 3.125 1.960 ;
        RECT  2.895 1.200 3.125 2.825 ;
        RECT  6.780 1.840 7.120 2.825 ;
        RECT  2.895 2.595 7.120 2.825 ;
        RECT  3.780 2.595 4.120 3.395 ;
        RECT  5.630 1.105 5.970 1.610 ;
        RECT  5.630 1.380 7.735 1.610 ;
        RECT  7.450 1.380 7.735 3.285 ;
        RECT  6.350 3.055 7.735 3.285 ;
        RECT  6.350 3.055 6.690 3.385 ;
    END
END HA1_X8_18_SVT_WB

MACRO HA1_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN HA1_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.940 2.165 5.090 2.395 ;
        RECT  4.570 1.820 5.090 2.395 ;
        RECT  1.940 1.860 2.280 2.395 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.800 1.620 4.080 1.935 ;
        RECT  2.800 1.260 3.270 1.935 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 2.330 1.240 3.135 ;
        RECT  0.900 0.685 1.240 1.385 ;
        RECT  0.700 1.045 0.930 2.710 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.605 1.675 7.140 3.280 ;
        RECT  6.605 0.535 6.900 3.280 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  7.370 2.470 7.660 4.100 ;
        RECT  5.800 3.545 6.140 4.100 ;
        RECT  3.140 3.110 4.180 4.100 ;
        RECT  1.700 3.110 2.040 4.100 ;
        RECT  0.180 2.600 0.470 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  7.280 -0.180 7.620 1.290 ;
        RECT  5.800 -0.180 6.140 0.820 ;
        RECT  1.660 -0.180 2.000 0.980 ;
        RECT  0.180 -0.180 0.470 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.550 0.535 5.330 0.875 ;
        RECT  3.550 0.535 3.890 1.280 ;
        RECT  2.340 0.745 3.190 1.030 ;
        RECT  2.340 0.745 2.570 1.550 ;
        RECT  1.470 1.210 2.570 1.550 ;
        RECT  1.160 1.620 1.700 1.960 ;
        RECT  1.470 1.210 1.700 2.855 ;
        RECT  5.420 1.840 5.760 2.855 ;
        RECT  1.470 2.625 5.760 2.855 ;
        RECT  2.420 2.625 2.760 3.395 ;
        RECT  4.270 1.105 4.610 1.480 ;
        RECT  4.270 1.250 6.375 1.480 ;
        RECT  6.090 1.250 6.375 3.315 ;
        RECT  4.990 3.085 6.375 3.315 ;
        RECT  4.990 3.085 5.330 3.385 ;
    END
END HA1_X4_18_SVT_WB

MACRO HA1_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN HA1_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.820 4.110 2.100 ;
        RECT  1.460 1.820 1.800 2.655 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.140 2.270 1.590 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.630 0.520 3.240 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.695 0.580 6.020 3.190 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  3.045 3.515 4.745 4.100 ;
        RECT  0.940 3.525 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.880 -0.180 5.220 0.405 ;
        RECT  0.940 -0.180 1.280 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.830 0.545 4.610 0.775 ;
        RECT  4.270 0.545 4.610 1.130 ;
        RECT  2.830 0.545 3.170 1.185 ;
        RECT  0.750 0.580 2.470 0.910 ;
        RECT  4.490 1.860 4.775 2.560 ;
        RECT  2.170 2.330 4.775 2.560 ;
        RECT  0.750 0.580 1.035 3.295 ;
        RECT  2.170 2.330 2.510 3.295 ;
        RECT  0.750 2.955 2.510 3.295 ;
        RECT  3.550 1.005 3.890 1.590 ;
        RECT  3.550 1.360 5.235 1.590 ;
        RECT  5.005 1.620 5.465 1.960 ;
        RECT  5.005 1.360 5.235 3.090 ;
        RECT  3.990 2.790 5.235 3.090 ;
    END
END HA1_X2_18_SVT_WB

MACRO HA1_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN HA1_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.795 4.060 2.135 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 1.095 2.505 1.560 ;
        END
    END B
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.640 0.760 0.980 ;
        RECT  0.245 0.640 0.530 3.450 ;
        RECT  0.140 0.640 0.530 1.335 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.435 2.930 6.020 3.270 ;
        RECT  5.710 0.805 6.020 3.270 ;
        RECT  5.480 0.805 6.020 1.105 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  3.925 3.515 4.220 4.100 ;
        RECT  3.465 3.515 3.695 4.100 ;
        RECT  2.940 3.515 3.235 4.100 ;
        RECT  1.005 3.010 1.290 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.880 -0.180 5.220 0.405 ;
        RECT  0.750 -0.180 1.090 0.365 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.780 0.410 4.560 0.640 ;
        RECT  4.220 0.410 4.560 1.105 ;
        RECT  2.780 0.410 3.120 1.155 ;
        RECT  1.010 0.595 2.280 0.865 ;
        RECT  1.010 0.595 1.290 2.705 ;
        RECT  4.420 2.255 4.745 2.595 ;
        RECT  0.760 2.365 4.745 2.595 ;
        RECT  0.760 2.365 2.520 2.705 ;
        RECT  1.765 2.365 2.520 3.450 ;
        RECT  3.500 0.870 3.840 1.565 ;
        RECT  3.500 1.335 5.480 1.565 ;
        RECT  4.245 1.335 5.480 1.650 ;
        RECT  4.975 1.335 5.480 1.675 ;
        RECT  4.975 1.335 5.205 3.115 ;
        RECT  3.940 2.825 5.205 3.115 ;
    END
END HA1_X1_18_SVT_WB

MACRO FILLTIE_18_SVT_WB
    CLASS CORE SPACER ;
    FOREIGN FILLTIE_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  0.540 2.970 0.880 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  0.540 -0.180 0.880 0.880 ;
        END
    END VSS
END FILLTIE_18_SVT_WB

MACRO FILLER_X8_18_SVT_WB
    CLASS CORE SPACER ;
    FOREIGN FILLER_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  0.165 3.570 4.315 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  0.180 -0.180 4.310 0.350 ;
        END
    END VSS
END FILLER_X8_18_SVT_WB

MACRO FILLER_X4_18_SVT_WB
    CLASS CORE SPACER ;
    FOREIGN FILLER_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.170 3.570 2.070 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.170 -0.180 2.075 0.350 ;
        END
    END VSS
END FILLER_X4_18_SVT_WB

MACRO FILLER_X32_18_SVT_WB
    CLASS CORE SPACER ;
    FOREIGN FILLER_X32_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.920 4.100 ;
        RECT  0.165 3.570 17.760 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.920 0.180 ;
        RECT  0.165 -0.180 17.755 0.350 ;
        END
    END VSS
END FILLER_X32_18_SVT_WB

MACRO FILLER_X2_18_SVT_WB
    CLASS CORE SPACER ;
    FOREIGN FILLER_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.120 4.100 ;
        RECT  0.400 3.570 0.740 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.120 0.180 ;
        RECT  0.370 -0.180 0.710 0.350 ;
        END
    END VSS
END FILLER_X2_18_SVT_WB

MACRO FILLER_X1_18_SVT_WB
    CLASS CORE SPACER ;
    FOREIGN FILLER_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 0.560 0.180 ;
        END
    END VSS
END FILLER_X1_18_SVT_WB

MACRO FILLER_X16_18_SVT_WB
    CLASS CORE SPACER ;
    FOREIGN FILLER_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  0.180 3.570 8.775 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  0.180 -0.180 8.755 0.350 ;
        END
    END VSS
END FILLER_X16_18_SVT_WB

MACRO FILLCAP_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN FILLCAP_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.120 2.380 3.460 4.100 ;
        RECT  2.400 2.380 2.740 4.100 ;
        RECT  0.960 2.375 1.300 4.100 ;
        RECT  0.240 2.430 0.580 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  2.680 -0.180 3.020 0.810 ;
        RECT  1.960 -0.180 2.300 0.810 ;
        RECT  1.240 -0.180 1.580 0.820 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.680 1.620 3.680 1.960 ;
        RECT  1.680 1.620 2.020 3.445 ;
        RECT  0.520 0.580 0.860 1.390 ;
        RECT  3.400 0.580 3.740 1.390 ;
        RECT  0.520 1.085 3.740 1.390 ;
        RECT  0.520 0.580 0.750 2.200 ;
        RECT  0.300 1.860 0.750 2.200 ;
    END
END FILLCAP_X8_18_SVT_WB

MACRO FILLCAP_X64_18_SVT_WB
    CLASS CORE ;
    FOREIGN FILLCAP_X64_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 25.760 4.100 ;
        RECT  23.420 2.600 23.760 4.100 ;
        RECT  22.700 2.600 23.040 4.100 ;
        RECT  21.260 2.600 21.600 4.100 ;
        RECT  20.540 2.600 20.880 4.100 ;
        RECT  19.820 2.600 20.160 4.100 ;
        RECT  18.380 2.600 18.720 4.100 ;
        RECT  17.660 2.600 18.000 4.100 ;
        RECT  16.940 2.600 17.280 4.100 ;
        RECT  15.500 2.600 15.840 4.100 ;
        RECT  14.780 2.600 15.120 4.100 ;
        RECT  14.060 2.600 14.400 4.100 ;
        RECT  12.620 2.600 12.960 4.100 ;
        RECT  11.900 2.595 12.240 4.100 ;
        RECT  11.180 2.595 11.520 4.100 ;
        RECT  9.740 2.595 10.080 4.100 ;
        RECT  9.020 2.595 9.360 4.100 ;
        RECT  8.300 2.640 8.640 4.100 ;
        RECT  6.860 2.435 7.200 4.100 ;
        RECT  6.140 2.600 6.480 4.100 ;
        RECT  5.420 2.600 5.760 4.100 ;
        RECT  3.980 2.600 4.320 4.100 ;
        RECT  3.260 2.600 3.600 4.100 ;
        RECT  2.540 3.110 2.880 4.100 ;
        RECT  1.100 2.445 1.440 4.100 ;
        RECT  0.380 2.445 0.720 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 25.760 0.180 ;
        RECT  24.120 -0.180 24.460 0.855 ;
        RECT  23.400 -0.180 23.740 0.810 ;
        RECT  22.680 -0.180 23.020 0.855 ;
        RECT  21.240 -0.180 21.580 0.855 ;
        RECT  20.520 -0.180 20.860 0.810 ;
        RECT  19.800 -0.180 20.140 0.855 ;
        RECT  18.360 -0.180 18.700 0.855 ;
        RECT  17.640 -0.180 17.980 0.810 ;
        RECT  16.920 -0.180 17.260 0.855 ;
        RECT  15.480 -0.180 15.820 0.855 ;
        RECT  14.760 -0.180 15.100 0.810 ;
        RECT  14.040 -0.180 14.380 0.810 ;
        RECT  12.600 -0.180 12.940 0.855 ;
        RECT  11.880 -0.180 12.220 0.810 ;
        RECT  11.160 -0.180 11.500 0.855 ;
        RECT  9.720 -0.180 10.060 0.855 ;
        RECT  9.000 -0.180 9.340 0.810 ;
        RECT  8.280 -0.180 8.620 0.855 ;
        RECT  6.840 -0.180 7.180 0.855 ;
        RECT  6.120 -0.180 6.460 0.810 ;
        RECT  5.400 -0.180 5.740 0.855 ;
        RECT  3.960 -0.180 4.300 0.855 ;
        RECT  3.240 -0.180 3.580 0.810 ;
        RECT  2.520 -0.180 2.860 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  4.680 0.515 5.020 1.325 ;
        RECT  7.560 0.515 7.900 1.325 ;
        RECT  10.440 0.515 10.780 1.325 ;
        RECT  13.320 0.515 13.660 1.325 ;
        RECT  16.200 0.515 16.540 1.325 ;
        RECT  19.080 0.515 19.420 1.325 ;
        RECT  21.960 0.515 22.300 1.325 ;
        RECT  24.840 0.515 25.180 1.325 ;
        RECT  1.800 1.085 25.180 1.325 ;
        RECT  1.800 0.470 2.140 2.200 ;
        RECT  0.200 1.860 2.140 2.200 ;
        RECT  2.370 1.620 25.400 1.960 ;
        RECT  2.370 1.620 2.710 2.775 ;
        RECT  1.820 2.435 2.710 2.775 ;
        RECT  4.700 1.620 5.040 3.190 ;
        RECT  13.340 1.620 13.680 3.190 ;
        RECT  16.220 1.620 16.560 3.190 ;
        RECT  19.100 1.620 19.440 3.190 ;
        RECT  21.980 1.620 22.320 3.190 ;
        RECT  1.820 2.435 2.160 3.245 ;
        RECT  7.580 1.620 7.920 3.245 ;
        RECT  10.460 1.620 10.800 3.405 ;
    END
END FILLCAP_X64_18_SVT_WB

MACRO FILLCAP_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN FILLCAP_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.230 2.430 0.570 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.670 -0.180 2.010 1.390 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.350 0.475 0.690 2.200 ;
        RECT  0.165 1.860 0.690 2.200 ;
        RECT  1.580 1.620 2.075 1.960 ;
        RECT  1.580 1.620 1.890 3.445 ;
    END
END FILLCAP_X4_18_SVT_WB

MACRO FILLCAP_X32_18_SVT_WB
    CLASS CORE ;
    FOREIGN FILLCAP_X32_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 13.440 4.100 ;
        RECT  11.750 2.625 12.090 4.100 ;
        RECT  11.005 2.600 11.405 4.100 ;
        RECT  9.590 2.625 9.930 4.100 ;
        RECT  8.865 2.600 9.235 4.100 ;
        RECT  8.150 2.625 8.490 4.100 ;
        RECT  6.710 2.625 7.050 4.100 ;
        RECT  5.975 2.630 6.350 4.100 ;
        RECT  5.270 2.635 5.610 4.100 ;
        RECT  3.830 2.635 4.170 4.100 ;
        RECT  3.110 2.620 3.455 4.100 ;
        RECT  2.390 2.635 2.730 4.100 ;
        RECT  0.935 2.620 1.305 4.100 ;
        RECT  0.230 2.645 0.570 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 13.440 0.180 ;
        RECT  12.190 -0.180 12.530 0.855 ;
        RECT  11.445 -0.180 11.845 0.855 ;
        RECT  10.750 -0.180 11.090 0.855 ;
        RECT  9.310 -0.180 9.650 0.855 ;
        RECT  8.590 -0.180 8.940 0.855 ;
        RECT  7.870 -0.180 8.210 0.855 ;
        RECT  6.430 -0.180 6.770 0.855 ;
        RECT  5.685 -0.180 6.065 0.855 ;
        RECT  4.990 -0.180 5.330 0.855 ;
        RECT  3.550 -0.180 3.890 0.855 ;
        RECT  2.810 -0.180 3.185 0.855 ;
        RECT  2.110 -0.180 2.450 0.855 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.700 1.620 13.250 1.960 ;
        RECT  7.430 1.620 7.770 3.215 ;
        RECT  1.700 1.620 2.010 3.225 ;
        RECT  10.310 1.620 10.650 3.230 ;
        RECT  4.550 1.620 4.890 3.235 ;
        RECT  1.390 0.515 1.730 1.325 ;
        RECT  4.270 0.515 4.610 1.325 ;
        RECT  7.150 0.515 7.490 1.325 ;
        RECT  10.030 0.515 10.370 1.325 ;
        RECT  12.910 0.515 13.250 1.325 ;
        RECT  1.240 1.085 13.250 1.325 ;
        RECT  1.240 1.050 1.470 2.195 ;
        RECT  0.245 1.855 1.470 2.195 ;
    END
END FILLCAP_X32_18_SVT_WB

MACRO FILLCAP_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN FILLCAP_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  5.940 2.380 6.280 4.100 ;
        RECT  5.190 2.570 5.575 4.100 ;
        RECT  3.780 2.595 4.120 4.100 ;
        RECT  2.340 2.600 2.680 4.100 ;
        RECT  0.895 2.380 1.240 4.100 ;
        RECT  0.180 2.430 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  5.480 -0.180 5.820 0.920 ;
        RECT  4.745 -0.180 5.110 0.840 ;
        RECT  4.040 -0.180 4.380 0.855 ;
        RECT  2.600 -0.180 2.940 0.855 ;
        RECT  1.880 -0.180 2.220 0.855 ;
        RECT  1.160 -0.180 1.500 0.855 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.620 1.620 6.500 1.960 ;
        RECT  1.620 1.620 1.960 3.190 ;
        RECT  4.500 1.620 4.840 3.410 ;
        RECT  0.440 0.580 0.780 1.390 ;
        RECT  3.320 0.515 3.660 1.390 ;
        RECT  0.440 1.085 3.660 1.390 ;
        RECT  6.200 0.580 6.540 1.390 ;
        RECT  0.440 1.150 6.540 1.390 ;
        RECT  0.440 0.580 0.670 2.200 ;
        RECT  0.220 1.860 0.670 2.200 ;
    END
END FILLCAP_X16_18_SVT_WB

MACRO FA1_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN FA1_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.145 1.200 3.890 1.545 ;
        RECT  3.145 1.200 3.585 1.905 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.890 1.995 4.360 2.715 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.591  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.170 1.535 10.580 1.875 ;
        RECT  4.590 1.535 10.580 1.775 ;
        RECT  4.590 1.535 5.160 2.345 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.040 2.310 14.380 3.390 ;
        RECT  12.720 1.045 14.380 1.385 ;
        RECT  14.040 0.575 14.380 1.385 ;
        RECT  13.405 1.045 14.050 2.670 ;
        RECT  12.720 2.320 14.380 2.670 ;
        RECT  12.720 2.320 13.060 3.385 ;
        RECT  12.720 0.580 13.060 1.385 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.075 2.540 2.370 3.445 ;
        RECT  0.755 0.950 2.370 1.345 ;
        RECT  2.075 0.485 2.370 1.345 ;
        RECT  0.755 2.540 2.370 2.880 ;
        RECT  1.085 0.950 1.745 2.880 ;
        RECT  0.755 2.540 1.095 3.445 ;
        RECT  0.755 0.485 1.095 1.345 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.120 4.100 ;
        RECT  11.960 3.515 12.300 4.100 ;
        RECT  9.290 3.025 9.630 4.100 ;
        RECT  7.870 2.565 8.210 4.100 ;
        RECT  6.390 3.035 6.730 4.100 ;
        RECT  2.835 3.515 3.175 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.120 0.180 ;
        RECT  12.000 -0.180 12.340 1.390 ;
        RECT  9.330 -0.180 9.670 0.845 ;
        RECT  7.870 -0.180 8.210 1.240 ;
        RECT  6.390 -0.180 6.730 0.845 ;
        RECT  2.835 -0.180 3.175 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.600 0.635 5.250 0.865 ;
        RECT  4.910 0.635 5.250 1.260 ;
        RECT  2.600 0.635 2.885 3.285 ;
        RECT  4.910 2.580 5.250 3.285 ;
        RECT  2.600 3.055 5.250 3.285 ;
        RECT  5.630 2.565 7.490 2.805 ;
        RECT  5.630 2.565 5.970 2.905 ;
        RECT  7.150 2.565 7.490 2.905 ;
        RECT  5.630 0.920 5.970 1.305 ;
        RECT  7.150 0.920 7.490 1.305 ;
        RECT  5.630 1.075 7.490 1.305 ;
        RECT  8.570 2.565 10.430 2.795 ;
        RECT  10.090 2.565 10.430 2.850 ;
        RECT  8.570 2.565 8.910 3.100 ;
        RECT  8.570 1.000 8.910 1.305 ;
        RECT  10.090 1.000 10.430 1.305 ;
        RECT  8.570 1.075 10.430 1.305 ;
        RECT  10.810 1.620 12.580 1.960 ;
        RECT  5.390 2.005 5.730 2.335 ;
        RECT  5.390 2.105 11.150 2.335 ;
        RECT  10.810 1.015 11.150 2.720 ;
    END
END FA1_X8_18_SVT_WB

MACRO FA1_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN FA1_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.210 2.235 1.780 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 2.320 2.860 2.660 ;
        RECT  2.520 2.005 2.860 2.660 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.591  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.505 1.535 9.100 1.875 ;
        RECT  3.210 1.535 9.100 1.765 ;
        RECT  3.210 1.535 3.780 2.290 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.255 0.575 11.620 3.385 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 0.535 1.050 3.385 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  10.480 3.515 10.820 4.100 ;
        RECT  7.810 3.025 8.150 4.100 ;
        RECT  6.390 2.565 6.730 4.100 ;
        RECT  4.910 3.035 5.250 4.100 ;
        RECT  1.515 3.515 1.855 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  10.520 -0.180 10.860 1.385 ;
        RECT  7.850 -0.180 8.190 0.845 ;
        RECT  6.390 -0.180 6.730 1.240 ;
        RECT  4.910 -0.180 5.250 0.845 ;
        RECT  1.515 -0.180 1.855 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.280 0.750 3.770 0.980 ;
        RECT  3.430 0.750 3.770 1.240 ;
        RECT  1.280 0.750 1.565 3.120 ;
        RECT  3.430 2.680 3.770 3.120 ;
        RECT  1.280 2.890 3.770 3.120 ;
        RECT  4.150 2.565 6.010 2.805 ;
        RECT  4.150 2.565 4.490 2.905 ;
        RECT  5.670 2.565 6.010 2.905 ;
        RECT  4.150 0.920 4.490 1.305 ;
        RECT  5.670 0.920 6.010 1.305 ;
        RECT  4.150 1.075 6.010 1.305 ;
        RECT  7.090 2.565 8.950 2.795 ;
        RECT  8.610 2.565 8.950 2.850 ;
        RECT  7.090 2.565 7.430 3.100 ;
        RECT  7.090 1.000 7.430 1.305 ;
        RECT  8.610 1.000 8.950 1.305 ;
        RECT  7.090 1.075 8.950 1.305 ;
        RECT  9.330 1.620 11.025 1.960 ;
        RECT  4.010 1.995 4.295 2.335 ;
        RECT  4.010 2.105 9.670 2.335 ;
        RECT  9.330 1.015 9.670 2.720 ;
    END
END FA1_X4_18_SVT_WB

MACRO FA1_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN FA1_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.210 1.675 1.780 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.560 2.305 2.300 2.660 ;
        RECT  1.960 2.005 2.300 2.660 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.548  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.955 1.535 8.555 1.875 ;
        RECT  2.650 1.535 8.555 1.765 ;
        RECT  2.650 1.535 3.220 2.235 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.520 2.590 11.060 3.290 ;
        RECT  10.680 0.530 11.060 3.290 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.550 0.490 3.385 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  9.760 3.515 10.100 4.100 ;
        RECT  7.250 3.035 7.590 4.100 ;
        RECT  5.830 2.605 6.170 4.100 ;
        RECT  4.350 3.025 4.690 4.100 ;
        RECT  0.945 3.515 1.285 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  9.920 -0.180 10.260 1.285 ;
        RECT  7.290 -0.180 7.630 0.845 ;
        RECT  5.830 -0.180 6.170 1.240 ;
        RECT  4.350 -0.180 4.690 0.845 ;
        RECT  0.945 -0.180 1.285 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.720 0.750 3.210 0.980 ;
        RECT  2.870 0.750 3.210 1.245 ;
        RECT  0.720 0.750 1.005 3.120 ;
        RECT  2.870 2.525 3.210 3.120 ;
        RECT  0.720 2.890 3.210 3.120 ;
        RECT  3.590 2.565 5.450 2.795 ;
        RECT  3.590 2.565 3.930 2.895 ;
        RECT  5.110 2.565 5.450 2.895 ;
        RECT  3.590 0.920 3.930 1.305 ;
        RECT  5.110 0.920 5.450 1.305 ;
        RECT  3.590 1.075 5.450 1.305 ;
        RECT  6.530 2.565 8.390 2.805 ;
        RECT  6.530 2.565 6.870 3.165 ;
        RECT  6.530 1.000 6.870 1.305 ;
        RECT  8.050 1.000 8.390 1.305 ;
        RECT  6.530 1.075 8.390 1.305 ;
        RECT  8.785 1.620 10.450 1.960 ;
        RECT  3.450 1.995 3.735 2.335 ;
        RECT  3.450 2.105 9.110 2.335 ;
        RECT  8.785 1.000 9.110 2.720 ;
        RECT  8.770 2.105 9.110 2.720 ;
    END
END FA1_X2_18_SVT_WB

MACRO FA1_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN FA1_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.605  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.330 2.545 9.465 2.875 ;
        RECT  9.100 2.100 9.465 2.875 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.605  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.760 1.975 8.830 2.315 ;
        RECT  8.490 1.615 8.830 2.315 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.505 8.130 1.745 ;
        RECT  2.380 1.045 2.770 1.745 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.155 0.805 10.500 2.960 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.890 0.480 3.030 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.560 3.565 10.370 4.100 ;
        RECT  5.530 3.110 5.870 4.100 ;
        RECT  0.340 3.565 1.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.615 -0.180 10.315 0.405 ;
        RECT  5.530 -0.180 5.870 0.810 ;
        RECT  0.270 -0.180 1.080 0.355 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.670 0.470 3.010 0.815 ;
        RECT  0.710 0.585 3.010 0.815 ;
        RECT  0.710 0.585 1.000 3.335 ;
        RECT  0.710 3.105 3.010 3.335 ;
        RECT  2.670 3.105 3.010 3.450 ;
        RECT  3.390 3.110 5.150 3.450 ;
        RECT  3.390 0.470 5.150 0.810 ;
        RECT  6.230 3.105 7.890 3.435 ;
        RECT  6.230 0.485 7.890 0.815 ;
        RECT  8.270 0.485 8.610 1.275 ;
        RECT  3.150 1.045 9.925 1.275 ;
        RECT  9.695 1.045 9.925 3.335 ;
        RECT  8.270 3.105 9.925 3.335 ;
        RECT  8.270 3.105 8.610 3.435 ;
    END
END FA1_X1_18_SVT_WB

MACRO FA1_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN FA1_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.605  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.575 9.950 2.815 ;
        RECT  9.610 2.475 9.950 2.815 ;
        RECT  1.210 2.380 1.590 2.815 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.605  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.890 2.095 9.380 2.345 ;
        RECT  8.940 1.770 9.380 2.345 ;
        RECT  1.890 2.005 2.190 2.345 ;
        END
    END B
    PIN CI
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.570 8.560 1.865 ;
        RECT  2.380 1.525 2.940 1.865 ;
        RECT  2.380 1.210 2.660 1.865 ;
        END
    END CI
    PIN CO
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.650 0.535 11.060 3.450 ;
        END
    END CO
    PIN S
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 0.535 0.465 3.385 ;
        END
    END S
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  9.890 3.515 10.230 4.100 ;
        RECT  7.220 3.515 7.560 4.100 ;
        RECT  5.760 3.045 6.100 4.100 ;
        RECT  4.280 3.515 4.620 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  9.890 -0.180 10.230 0.875 ;
        RECT  7.220 -0.180 7.560 0.405 ;
        RECT  5.760 -0.180 6.100 0.875 ;
        RECT  4.280 -0.180 4.620 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.800 0.535 3.140 0.915 ;
        RECT  0.695 0.685 3.140 0.915 ;
        RECT  0.695 0.685 0.980 3.285 ;
        RECT  0.695 3.045 3.140 3.285 ;
        RECT  2.800 3.045 3.140 3.385 ;
        RECT  3.520 3.045 5.380 3.285 ;
        RECT  3.520 3.045 3.860 3.385 ;
        RECT  5.040 3.045 5.380 3.385 ;
        RECT  3.520 0.535 3.860 0.875 ;
        RECT  5.040 0.535 5.380 0.875 ;
        RECT  3.520 0.635 5.380 0.875 ;
        RECT  6.460 3.045 8.320 3.285 ;
        RECT  6.460 3.045 6.800 3.385 ;
        RECT  7.980 3.045 8.320 3.385 ;
        RECT  6.460 0.535 6.800 0.875 ;
        RECT  7.980 0.535 8.320 0.875 ;
        RECT  6.460 0.635 8.320 0.875 ;
        RECT  8.700 0.535 9.040 1.340 ;
        RECT  3.280 1.105 10.420 1.340 ;
        RECT  8.910 1.105 10.420 1.445 ;
        RECT  10.180 1.105 10.420 3.285 ;
        RECT  8.700 3.045 10.420 3.285 ;
        RECT  8.700 3.045 9.040 3.385 ;
    END
END FA1_X0_18_SVT_WB

MACRO DLY4_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY4_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.756  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.735 0.825 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.254  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.770 0.535 3.250 3.415 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.460 3.080 2.360 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  1.500 -0.180 2.320 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.460 1.720 2.280 2.060 ;
        RECT  1.460 1.100 1.800 2.720 ;
    END
END DLY4_X4_18_SVT_WB

MACRO DLY4_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY4_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.756  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.735 0.945 2.280 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.526  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.735 0.535 3.245 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.460 3.080 2.355 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.500 -0.180 2.315 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.460 1.720 2.275 2.060 ;
        RECT  1.460 1.100 1.800 2.720 ;
    END
END DLY4_X1_18_SVT_WB

MACRO DLY3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.605  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.735 0.825 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.364  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.640 0.535 3.225 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.455 2.370 3.765 4.100 ;
        RECT  1.280 3.080 2.180 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.455 -0.180 3.735 1.465 ;
        RECT  1.320 -0.180 2.140 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.280 1.720 2.100 2.060 ;
        RECT  1.280 1.100 1.620 2.720 ;
    END
END DLY3_X4_18_SVT_WB

MACRO DLY3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.605  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.200 1.735 1.005 2.280 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.526  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.710 0.535 3.240 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.340 3.080 2.330 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.380 -0.180 2.290 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.340 1.720 2.250 2.060 ;
        RECT  1.340 1.100 1.680 2.720 ;
    END
END DLY3_X1_18_SVT_WB

MACRO DLY2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.300 1.735 1.005 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.364  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.640 0.535 3.225 3.365 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  3.455 2.365 3.760 4.100 ;
        RECT  1.280 3.080 2.180 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.455 -0.180 3.750 1.430 ;
        RECT  1.320 -0.180 2.140 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.280 1.720 2.100 2.060 ;
        RECT  1.280 1.100 1.620 2.720 ;
    END
END DLY2_X4_18_SVT_WB

MACRO DLY2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.240 1.735 1.005 2.280 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.526  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.710 0.535 3.240 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.340 3.080 2.330 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.380 -0.180 2.290 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.340 1.720 2.250 2.060 ;
        RECT  1.340 1.100 1.680 2.720 ;
    END
END DLY2_X1_18_SVT_WB

MACRO DLY1_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY1_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.735 0.710 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.535 2.690 3.355 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.940 3.080 1.830 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.980 -0.180 1.790 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 1.720 1.750 2.060 ;
        RECT  0.940 1.100 1.280 2.720 ;
    END
END DLY1_X4_18_SVT_WB

MACRO DLY1_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DLY1_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.735 0.710 2.220 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.526  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.210 0.535 2.660 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.940 3.080 1.830 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.980 -0.180 1.790 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 1.720 1.750 2.060 ;
        RECT  0.940 1.100 1.280 2.720 ;
    END
END DLY1_X1_18_SVT_WB

MACRO DFF_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFF_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.530 0.760 2.295 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.211  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.450 3.295 2.110 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.680 0.535 11.060 3.385 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.172  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.155 1.105 8.385 2.705 ;
        RECT  7.945 2.430 8.230 3.385 ;
        RECT  7.880 1.105 8.385 1.540 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  9.920 3.515 10.260 4.100 ;
        RECT  7.120 3.540 7.460 4.100 ;
        RECT  4.505 2.550 4.845 4.100 ;
        RECT  2.100 2.415 2.440 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  9.920 -0.180 10.260 0.405 ;
        RECT  7.120 -0.180 7.460 0.405 ;
        RECT  2.200 -0.180 2.540 0.350 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.945 0.520 1.300 ;
        RECT  0.180 1.070 1.375 1.300 ;
        RECT  1.090 1.070 1.375 2.865 ;
        RECT  0.180 2.525 1.375 2.865 ;
        RECT  3.250 0.880 4.915 1.220 ;
        RECT  4.630 0.880 4.915 1.860 ;
        RECT  3.525 0.880 3.755 2.790 ;
        RECT  3.250 2.450 3.755 2.790 ;
        RECT  3.985 1.980 4.300 2.320 ;
        RECT  5.145 1.000 5.580 2.320 ;
        RECT  3.985 2.090 5.580 2.320 ;
        RECT  5.265 1.000 5.580 3.090 ;
        RECT  2.765 0.410 6.640 0.650 ;
        RECT  1.500 0.580 2.990 0.875 ;
        RECT  1.640 0.580 2.100 2.185 ;
        RECT  6.380 0.410 6.640 2.570 ;
        RECT  6.300 2.230 6.640 2.570 ;
        RECT  1.640 0.580 1.870 3.390 ;
        RECT  1.515 3.050 1.870 3.390 ;
        RECT  5.810 0.880 6.150 1.220 ;
        RECT  7.485 1.860 7.925 2.200 ;
        RECT  5.810 0.880 6.070 3.310 ;
        RECT  7.485 1.860 7.715 3.310 ;
        RECT  5.810 2.970 7.715 3.310 ;
        RECT  9.160 0.535 9.500 0.875 ;
        RECT  6.970 0.635 10.450 0.875 ;
        RECT  6.970 0.635 7.255 1.980 ;
        RECT  10.165 0.635 10.450 3.285 ;
        RECT  9.160 3.045 10.450 3.285 ;
        RECT  9.160 3.045 9.500 3.385 ;
    END
END DFF_X4_18_SVT_WB

MACRO DFF_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFF_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.525 0.745 2.285 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.211  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.485 3.445 2.170 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.982  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.120 0.470 10.500 3.380 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.032  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.255 1.100 8.485 2.770 ;
        RECT  8.035 2.430 8.320 3.385 ;
        RECT  7.930 1.100 8.485 1.540 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  9.400 3.040 9.740 4.100 ;
        RECT  7.220 3.515 7.560 4.100 ;
        RECT  4.630 2.545 4.970 4.100 ;
        RECT  2.250 2.565 2.590 4.100 ;
        RECT  0.740 3.510 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  9.400 -0.180 9.740 0.810 ;
        RECT  7.220 -0.180 7.560 0.400 ;
        RECT  2.290 -0.180 2.630 0.350 ;
        RECT  0.830 -0.180 1.170 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.955 0.520 1.295 ;
        RECT  0.180 1.060 1.430 1.295 ;
        RECT  1.090 1.060 1.430 2.810 ;
        RECT  0.180 2.515 1.430 2.810 ;
        RECT  3.400 0.915 5.160 1.255 ;
        RECT  4.870 0.915 5.160 1.815 ;
        RECT  3.675 0.915 3.905 2.755 ;
        RECT  3.400 2.415 3.905 2.755 ;
        RECT  4.135 1.945 4.450 2.285 ;
        RECT  4.135 2.045 5.730 2.285 ;
        RECT  5.390 0.915 5.730 3.105 ;
        RECT  2.855 0.410 6.830 0.685 ;
        RECT  1.590 0.580 3.080 0.890 ;
        RECT  1.730 0.580 2.120 2.235 ;
        RECT  6.600 0.410 6.830 2.585 ;
        RECT  6.445 2.245 6.830 2.585 ;
        RECT  1.730 0.580 1.960 3.380 ;
        RECT  1.500 3.040 1.960 3.380 ;
        RECT  5.985 0.915 6.370 1.255 ;
        RECT  7.575 1.860 8.025 2.200 ;
        RECT  5.985 0.915 6.215 3.225 ;
        RECT  7.575 1.860 7.805 3.225 ;
        RECT  5.985 2.885 7.805 3.225 ;
        RECT  7.060 0.630 9.020 0.870 ;
        RECT  7.060 0.630 7.345 1.980 ;
        RECT  8.715 1.640 9.890 1.980 ;
        RECT  8.715 0.630 9.020 3.240 ;
    END
END DFF_X2_18_SVT_WB

MACRO DFF_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFF_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.555 0.760 2.340 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.710 3.355 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.560 2.330 9.940 2.875 ;
        RECT  9.710 0.995 9.940 2.875 ;
        RECT  9.560 0.995 9.940 1.335 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.491  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.795 2.425 8.405 2.765 ;
        RECT  8.065 1.130 8.405 2.765 ;
        RECT  7.735 1.130 8.405 1.540 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  9.000 3.515 9.340 4.100 ;
        RECT  6.975 3.510 7.315 4.100 ;
        RECT  4.430 2.680 4.770 4.100 ;
        RECT  2.070 2.380 2.390 4.100 ;
        RECT  0.740 3.510 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  9.000 -0.180 9.340 0.410 ;
        RECT  6.975 -0.180 7.315 0.410 ;
        RECT  2.200 -0.180 2.540 0.350 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.985 0.520 1.325 ;
        RECT  0.180 1.060 1.375 1.325 ;
        RECT  1.090 1.060 1.375 2.855 ;
        RECT  0.180 2.570 1.375 2.855 ;
        RECT  3.215 0.880 4.920 1.220 ;
        RECT  4.580 0.880 4.920 1.740 ;
        RECT  3.630 0.880 3.970 2.770 ;
        RECT  3.200 2.430 3.970 2.770 ;
        RECT  4.205 2.110 5.490 2.450 ;
        RECT  5.150 0.880 5.490 3.020 ;
        RECT  2.765 0.410 6.615 0.650 ;
        RECT  1.500 0.580 2.985 0.865 ;
        RECT  1.610 0.580 2.100 2.150 ;
        RECT  6.385 0.410 6.615 2.515 ;
        RECT  6.205 2.175 6.615 2.515 ;
        RECT  1.610 0.580 1.840 3.390 ;
        RECT  1.500 3.050 1.840 3.390 ;
        RECT  5.745 0.880 6.155 1.220 ;
        RECT  7.335 1.870 7.835 2.195 ;
        RECT  5.745 0.880 5.975 3.070 ;
        RECT  7.335 1.870 7.565 3.070 ;
        RECT  5.745 2.745 7.565 3.070 ;
        RECT  8.215 0.430 8.555 0.870 ;
        RECT  6.845 0.640 9.330 0.870 ;
        RECT  9.100 1.555 9.480 1.895 ;
        RECT  6.845 0.640 7.105 1.990 ;
        RECT  9.100 0.640 9.330 3.285 ;
        RECT  8.240 3.055 9.330 3.285 ;
        RECT  8.240 3.055 8.580 3.465 ;
    END
END DFF_X1_18_SVT_WB

MACRO DFFTR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFTR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.595 0.795 2.325 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.915 1.775 3.520 2.200 ;
        RECT  2.915 1.495 3.320 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.885 0.470 12.430 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.050 2.480 9.695 2.775 ;
        RECT  9.465 1.145 9.695 2.775 ;
        RECT  9.050 1.145 9.695 1.570 ;
        RECT  9.050 2.480 9.430 3.255 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.255 1.495 2.685 2.200 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 13.440 4.100 ;
        RECT  12.805 2.665 13.215 4.100 ;
        RECT  11.310 3.110 11.650 4.100 ;
        RECT  8.430 3.485 8.770 4.100 ;
        RECT  5.915 2.700 6.255 4.100 ;
        RECT  2.935 2.950 3.275 4.100 ;
        RECT  0.740 3.370 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 13.440 0.180 ;
        RECT  12.800 -0.180 13.240 1.290 ;
        RECT  11.310 -0.180 11.650 0.810 ;
        RECT  8.430 -0.180 8.770 0.455 ;
        RECT  2.345 -0.180 2.685 0.365 ;
        RECT  0.810 -0.180 1.150 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.080 1.375 1.365 ;
        RECT  1.090 1.080 1.375 2.840 ;
        RECT  0.180 2.555 1.375 2.840 ;
        RECT  3.455 0.975 3.980 1.265 ;
        RECT  3.750 0.975 3.980 2.720 ;
        RECT  2.175 2.430 3.980 2.720 ;
        RECT  4.670 1.450 6.440 1.790 ;
        RECT  4.670 0.930 4.980 2.720 ;
        RECT  6.440 0.930 6.920 1.220 ;
        RECT  5.670 2.130 6.920 2.470 ;
        RECT  6.670 0.930 6.920 3.020 ;
        RECT  6.635 2.130 6.920 3.020 ;
        RECT  2.915 0.410 7.935 0.700 ;
        RECT  1.570 0.595 4.440 0.745 ;
        RECT  1.570 0.595 3.225 0.945 ;
        RECT  7.675 0.410 7.935 2.500 ;
        RECT  4.210 0.410 4.440 3.230 ;
        RECT  4.210 2.900 4.520 3.230 ;
        RECT  1.605 0.595 1.910 3.390 ;
        RECT  8.950 1.800 9.235 2.250 ;
        RECT  8.165 2.020 9.235 2.250 ;
        RECT  7.160 0.930 7.445 3.020 ;
        RECT  8.165 2.020 8.395 3.020 ;
        RECT  7.160 2.730 8.395 3.020 ;
        RECT  10.450 0.470 10.805 0.915 ;
        RECT  8.390 0.685 10.805 0.915 ;
        RECT  8.390 0.685 8.620 1.790 ;
        RECT  8.165 1.450 8.620 1.790 ;
        RECT  10.575 1.860 11.645 2.200 ;
        RECT  10.575 0.470 10.805 3.450 ;
        RECT  10.450 3.110 10.805 3.450 ;
    END
END DFFTR_X4_18_SVT_WB

MACRO DFFTR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFTR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.595 0.795 2.325 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.915 1.775 3.520 2.200 ;
        RECT  2.915 1.495 3.320 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.325 0.470 11.850 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.310 1.145 9.610 2.775 ;
        RECT  9.050 2.480 9.430 3.255 ;
        RECT  9.050 1.145 9.610 1.570 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.255 1.495 2.685 2.200 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  10.750 3.110 11.090 4.100 ;
        RECT  8.430 3.485 8.770 4.100 ;
        RECT  5.915 2.700 6.255 4.100 ;
        RECT  2.935 2.950 3.275 4.100 ;
        RECT  0.740 3.370 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  10.750 -0.180 11.090 0.810 ;
        RECT  8.430 -0.180 8.770 0.455 ;
        RECT  2.345 -0.180 2.685 0.365 ;
        RECT  0.810 -0.180 1.150 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.080 1.375 1.365 ;
        RECT  1.090 1.080 1.375 2.840 ;
        RECT  0.180 2.555 1.375 2.840 ;
        RECT  3.455 0.975 3.980 1.265 ;
        RECT  3.750 0.975 3.980 2.720 ;
        RECT  2.175 2.430 3.980 2.720 ;
        RECT  4.670 1.450 6.440 1.790 ;
        RECT  4.670 0.930 4.980 2.720 ;
        RECT  6.440 0.930 6.920 1.220 ;
        RECT  5.670 2.130 6.920 2.470 ;
        RECT  6.670 0.930 6.920 3.020 ;
        RECT  6.635 2.130 6.920 3.020 ;
        RECT  2.915 0.410 7.935 0.700 ;
        RECT  1.570 0.595 4.440 0.745 ;
        RECT  1.570 0.595 3.225 0.945 ;
        RECT  7.675 0.410 7.935 2.500 ;
        RECT  4.210 0.410 4.440 3.230 ;
        RECT  4.210 2.900 4.520 3.230 ;
        RECT  1.605 0.595 1.910 3.390 ;
        RECT  8.850 1.800 9.080 2.250 ;
        RECT  8.165 2.020 9.080 2.250 ;
        RECT  7.160 0.930 7.445 3.020 ;
        RECT  8.165 2.020 8.395 3.020 ;
        RECT  7.160 2.730 8.395 3.020 ;
        RECT  9.890 0.470 10.245 0.915 ;
        RECT  8.390 0.685 10.245 0.915 ;
        RECT  8.390 0.685 8.620 1.790 ;
        RECT  8.165 1.450 8.620 1.790 ;
        RECT  10.015 1.860 11.085 2.200 ;
        RECT  10.015 0.470 10.245 3.450 ;
        RECT  9.890 3.110 10.245 3.450 ;
    END
END DFFTR_X2_18_SVT_WB

MACRO DFFTR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFTR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.595 0.795 2.325 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.915 1.775 3.520 2.200 ;
        RECT  2.915 1.495 3.320 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.325 0.470 11.850 3.450 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.310 1.145 9.610 2.775 ;
        RECT  9.050 2.480 9.430 3.255 ;
        RECT  9.050 1.145 9.610 1.570 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.183  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.255 1.495 2.685 2.200 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  10.750 3.110 11.090 4.100 ;
        RECT  8.430 3.485 8.770 4.100 ;
        RECT  5.915 2.700 6.255 4.100 ;
        RECT  2.935 2.950 3.275 4.100 ;
        RECT  0.740 3.370 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  10.750 -0.180 11.090 0.810 ;
        RECT  8.430 -0.180 8.770 0.455 ;
        RECT  2.345 -0.180 2.685 0.365 ;
        RECT  0.810 -0.180 1.150 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.080 1.375 1.365 ;
        RECT  1.090 1.080 1.375 2.840 ;
        RECT  0.180 2.555 1.375 2.840 ;
        RECT  3.455 0.975 3.980 1.265 ;
        RECT  3.750 0.975 3.980 2.720 ;
        RECT  2.175 2.430 3.980 2.720 ;
        RECT  4.670 1.450 6.440 1.790 ;
        RECT  4.670 0.930 4.980 2.720 ;
        RECT  6.440 0.930 6.920 1.220 ;
        RECT  5.670 2.130 6.920 2.470 ;
        RECT  6.670 0.930 6.920 3.020 ;
        RECT  6.635 2.130 6.920 3.020 ;
        RECT  2.915 0.410 7.935 0.700 ;
        RECT  1.570 0.595 4.440 0.745 ;
        RECT  1.570 0.595 3.225 0.945 ;
        RECT  7.675 0.410 7.935 2.500 ;
        RECT  4.210 0.410 4.440 3.230 ;
        RECT  4.210 2.900 4.520 3.230 ;
        RECT  1.605 0.595 1.910 3.390 ;
        RECT  8.850 1.800 9.080 2.250 ;
        RECT  8.165 2.020 9.080 2.250 ;
        RECT  7.160 0.930 7.445 3.020 ;
        RECT  8.165 2.020 8.395 3.020 ;
        RECT  7.160 2.730 8.395 3.020 ;
        RECT  9.890 0.470 10.245 0.915 ;
        RECT  8.390 0.685 10.245 0.915 ;
        RECT  8.390 0.685 8.620 1.790 ;
        RECT  8.165 1.450 8.620 1.790 ;
        RECT  10.015 1.860 11.085 2.200 ;
        RECT  10.015 0.470 10.245 3.450 ;
        RECT  9.890 3.110 10.245 3.450 ;
    END
END DFFTR_X1_18_SVT_WB

MACRO DFFS_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFS_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.208  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.695 3.340 2.155 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.195 1.735 13.540 3.175 ;
        RECT  13.200 1.095 13.540 3.175 ;
        RECT  11.880 1.735 13.540 2.100 ;
        RECT  11.880 1.100 12.220 3.175 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.080 0.470 16.420 3.450 ;
        RECT  14.655 1.790 16.420 2.110 ;
        RECT  14.655 0.470 15.180 3.450 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.600 8.910 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.360 4.100 ;
        RECT  16.800 2.640 17.140 4.100 ;
        RECT  15.410 2.640 15.700 4.100 ;
        RECT  13.920 2.695 14.260 4.100 ;
        RECT  11.205 2.640 11.500 4.100 ;
        RECT  8.815 3.515 9.985 4.100 ;
        RECT  4.635 3.530 5.915 4.100 ;
        RECT  1.970 3.530 2.310 4.100 ;
        RECT  0.740 3.530 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.360 0.180 ;
        RECT  16.800 -0.180 17.140 1.275 ;
        RECT  15.410 -0.180 15.700 1.280 ;
        RECT  11.120 -0.180 11.460 0.405 ;
        RECT  9.460 -0.180 9.800 0.405 ;
        RECT  4.395 -0.180 4.735 0.365 ;
        RECT  2.100 -0.180 2.440 0.365 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.295 1.055 3.800 1.395 ;
        RECT  3.570 2.090 5.255 2.325 ;
        RECT  3.570 1.055 3.800 2.840 ;
        RECT  3.295 2.555 3.800 2.840 ;
        RECT  4.245 1.055 5.870 1.395 ;
        RECT  4.245 1.055 4.585 1.860 ;
        RECT  5.530 1.055 5.870 2.840 ;
        RECT  5.530 2.435 6.705 2.840 ;
        RECT  5.105 2.555 6.705 2.840 ;
        RECT  0.180 0.930 1.270 1.270 ;
        RECT  1.040 1.575 1.620 1.915 ;
        RECT  0.180 2.535 1.270 2.875 ;
        RECT  1.040 0.930 1.270 3.300 ;
        RECT  0.930 2.535 1.270 3.300 ;
        RECT  0.930 3.070 6.855 3.300 ;
        RECT  3.515 3.070 3.855 3.510 ;
        RECT  6.515 3.070 6.855 3.510 ;
        RECT  3.575 0.410 3.915 0.825 ;
        RECT  2.020 0.595 7.850 0.825 ;
        RECT  1.500 0.975 2.360 1.315 ;
        RECT  6.100 0.595 6.330 2.200 ;
        RECT  7.600 0.595 7.850 2.160 ;
        RECT  6.100 1.860 6.515 2.200 ;
        RECT  2.020 0.595 2.360 2.545 ;
        RECT  1.500 2.315 2.360 2.545 ;
        RECT  1.500 2.315 1.840 2.840 ;
        RECT  6.560 1.055 6.845 1.565 ;
        RECT  6.560 1.335 7.370 1.565 ;
        RECT  7.085 1.335 7.370 3.180 ;
        RECT  9.980 1.860 10.265 3.180 ;
        RECT  7.085 2.950 10.265 3.180 ;
        RECT  10.220 1.095 10.725 1.630 ;
        RECT  9.290 1.400 10.725 1.630 ;
        RECT  10.495 1.095 10.725 3.450 ;
        RECT  9.290 1.400 9.630 1.915 ;
        RECT  10.495 1.640 10.975 3.450 ;
        RECT  8.080 0.635 14.425 0.865 ;
        RECT  8.080 0.635 8.505 1.370 ;
        RECT  14.140 0.635 14.425 2.200 ;
        RECT  8.080 0.635 8.310 2.720 ;
        RECT  8.080 2.380 9.410 2.720 ;
        RECT  7.805 2.390 9.410 2.720 ;
    END
END DFFS_X8_18_SVT_WB

MACRO DFFS_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFS_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.208  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.770 3.340 2.230 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.880 1.100 12.220 3.145 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.335 0.470 13.860 3.450 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.218  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.600 8.910 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.560 4.100 ;
        RECT  14.090 2.640 14.380 4.100 ;
        RECT  12.600 2.695 12.940 4.100 ;
        RECT  8.505 3.515 10.165 4.100 ;
        RECT  9.825 3.465 10.165 4.100 ;
        RECT  4.635 3.530 5.915 4.100 ;
        RECT  2.105 3.530 2.445 4.100 ;
        RECT  0.740 3.530 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.560 0.180 ;
        RECT  14.090 -0.180 14.380 1.280 ;
        RECT  11.120 -0.180 11.460 0.405 ;
        RECT  9.535 -0.180 9.875 0.405 ;
        RECT  4.395 -0.180 4.735 0.365 ;
        RECT  2.100 -0.180 2.440 0.365 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.295 1.055 3.800 1.395 ;
        RECT  3.570 2.090 5.255 2.325 ;
        RECT  3.570 1.055 3.800 2.840 ;
        RECT  3.295 2.555 3.800 2.840 ;
        RECT  4.245 1.055 5.870 1.395 ;
        RECT  4.245 1.055 4.585 1.860 ;
        RECT  5.530 1.055 5.870 2.840 ;
        RECT  5.530 2.435 6.705 2.840 ;
        RECT  5.105 2.555 6.705 2.840 ;
        RECT  0.180 1.060 1.270 1.400 ;
        RECT  1.040 1.615 1.600 1.925 ;
        RECT  0.180 2.380 1.270 2.720 ;
        RECT  1.040 1.060 1.270 3.300 ;
        RECT  0.930 2.380 1.270 3.300 ;
        RECT  0.930 3.070 6.855 3.300 ;
        RECT  3.515 3.070 3.855 3.510 ;
        RECT  6.515 3.070 6.855 3.510 ;
        RECT  3.575 0.410 3.915 0.825 ;
        RECT  2.060 0.595 7.850 0.825 ;
        RECT  1.500 1.060 2.360 1.385 ;
        RECT  6.100 0.595 6.330 2.200 ;
        RECT  7.600 0.595 7.850 1.915 ;
        RECT  6.100 1.860 6.515 2.200 ;
        RECT  1.830 1.060 2.360 2.375 ;
        RECT  2.060 0.595 2.360 2.375 ;
        RECT  1.500 2.375 2.060 2.720 ;
        RECT  6.560 1.055 6.845 1.565 ;
        RECT  6.560 1.335 7.370 1.565 ;
        RECT  10.070 1.915 10.410 2.370 ;
        RECT  9.650 2.140 10.410 2.370 ;
        RECT  7.085 1.335 7.370 3.180 ;
        RECT  9.650 2.140 9.990 3.180 ;
        RECT  7.085 2.950 9.990 3.180 ;
        RECT  10.295 1.095 10.640 1.685 ;
        RECT  9.285 1.455 11.145 1.685 ;
        RECT  9.285 1.455 9.625 1.910 ;
        RECT  10.640 1.455 11.145 1.960 ;
        RECT  10.640 1.455 10.925 3.280 ;
        RECT  10.585 2.525 10.925 3.280 ;
        RECT  9.405 0.635 13.105 0.865 ;
        RECT  9.405 0.635 9.745 1.225 ;
        RECT  8.080 0.995 9.745 1.225 ;
        RECT  8.080 0.995 8.685 1.370 ;
        RECT  12.820 0.635 13.105 2.200 ;
        RECT  8.080 0.995 8.310 2.720 ;
        RECT  7.805 2.380 9.405 2.720 ;
    END
END DFFS_X4_18_SVT_WB

MACRO DFFS_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFS_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.208  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.770 3.340 2.230 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.320 1.100 11.690 3.205 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.000 0.525 13.300 2.855 ;
        RECT  12.750 2.490 13.105 3.400 ;
        RECT  12.775 0.525 13.300 1.450 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.218  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.600 8.910 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 13.440 4.100 ;
        RECT  12.040 3.020 12.380 4.100 ;
        RECT  8.505 3.515 10.165 4.100 ;
        RECT  9.825 3.465 10.165 4.100 ;
        RECT  4.635 3.530 5.915 4.100 ;
        RECT  2.105 3.530 2.445 4.100 ;
        RECT  0.740 3.530 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 13.440 0.180 ;
        RECT  9.535 -0.180 9.875 0.405 ;
        RECT  4.395 -0.180 4.735 0.365 ;
        RECT  2.100 -0.180 2.440 0.365 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.295 1.055 3.800 1.395 ;
        RECT  3.570 2.090 5.255 2.325 ;
        RECT  3.570 1.055 3.800 2.840 ;
        RECT  3.295 2.555 3.800 2.840 ;
        RECT  4.245 1.055 5.870 1.395 ;
        RECT  4.245 1.055 4.585 1.860 ;
        RECT  5.530 1.055 5.870 2.840 ;
        RECT  5.530 2.435 6.705 2.840 ;
        RECT  5.105 2.555 6.705 2.840 ;
        RECT  0.180 1.060 1.270 1.400 ;
        RECT  1.040 1.615 1.600 1.925 ;
        RECT  0.180 2.380 1.270 2.720 ;
        RECT  1.040 1.060 1.270 3.300 ;
        RECT  0.930 2.380 1.270 3.300 ;
        RECT  0.930 3.070 6.855 3.300 ;
        RECT  3.515 3.070 3.855 3.510 ;
        RECT  6.515 3.070 6.855 3.510 ;
        RECT  3.575 0.410 3.915 0.825 ;
        RECT  2.060 0.595 7.850 0.825 ;
        RECT  1.500 1.060 2.360 1.385 ;
        RECT  6.100 0.595 6.330 2.200 ;
        RECT  7.600 0.595 7.850 1.915 ;
        RECT  6.100 1.860 6.515 2.200 ;
        RECT  1.830 1.060 2.360 2.375 ;
        RECT  2.060 0.595 2.360 2.375 ;
        RECT  1.500 2.375 2.060 2.720 ;
        RECT  6.560 1.055 6.845 1.565 ;
        RECT  6.560 1.335 7.370 1.565 ;
        RECT  10.070 1.915 10.410 2.370 ;
        RECT  9.650 2.140 10.410 2.370 ;
        RECT  7.085 1.335 7.370 3.180 ;
        RECT  9.650 2.140 9.990 3.180 ;
        RECT  7.085 2.950 9.990 3.180 ;
        RECT  10.295 1.095 10.640 1.685 ;
        RECT  9.285 1.455 11.090 1.685 ;
        RECT  9.285 1.455 9.625 1.910 ;
        RECT  10.640 1.455 11.090 1.960 ;
        RECT  10.640 1.455 10.925 3.280 ;
        RECT  10.585 2.525 10.925 3.280 ;
        RECT  9.405 0.635 12.545 0.865 ;
        RECT  9.405 0.635 9.745 1.225 ;
        RECT  8.080 0.995 9.745 1.225 ;
        RECT  8.080 0.995 8.685 1.370 ;
        RECT  12.260 0.635 12.545 2.200 ;
        RECT  8.080 0.995 8.310 2.720 ;
        RECT  7.805 2.380 9.405 2.720 ;
    END
END DFFS_X2_18_SVT_WB

MACRO DFFS_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFS_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.208  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.770 3.340 2.230 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.320 1.100 11.690 2.745 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.775 2.490 13.300 2.855 ;
        RECT  13.000 1.035 13.300 2.855 ;
        RECT  12.775 1.035 13.300 1.450 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.218  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.600 8.910 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 13.440 4.100 ;
        RECT  8.505 3.515 10.165 4.100 ;
        RECT  9.825 3.465 10.165 4.100 ;
        RECT  4.635 3.530 5.915 4.100 ;
        RECT  2.105 3.530 2.445 4.100 ;
        RECT  0.740 3.530 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 13.440 0.180 ;
        RECT  9.535 -0.180 9.875 0.405 ;
        RECT  4.395 -0.180 4.735 0.365 ;
        RECT  2.100 -0.180 2.440 0.365 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.295 1.055 3.800 1.395 ;
        RECT  3.570 2.090 5.255 2.325 ;
        RECT  3.570 1.055 3.800 2.840 ;
        RECT  3.295 2.555 3.800 2.840 ;
        RECT  4.245 1.055 5.870 1.395 ;
        RECT  4.245 1.055 4.585 1.860 ;
        RECT  5.530 1.055 5.870 2.840 ;
        RECT  5.530 2.435 6.705 2.840 ;
        RECT  5.105 2.555 6.705 2.840 ;
        RECT  0.180 1.060 1.270 1.400 ;
        RECT  1.040 1.615 1.600 1.925 ;
        RECT  0.180 2.380 1.270 2.720 ;
        RECT  1.040 1.060 1.270 3.300 ;
        RECT  0.930 2.380 1.270 3.300 ;
        RECT  0.930 3.070 6.855 3.300 ;
        RECT  3.515 3.070 3.855 3.510 ;
        RECT  6.515 3.070 6.855 3.510 ;
        RECT  3.575 0.410 3.915 0.825 ;
        RECT  2.060 0.595 7.850 0.825 ;
        RECT  1.500 1.060 2.360 1.385 ;
        RECT  6.100 0.595 6.330 2.200 ;
        RECT  7.600 0.595 7.850 1.915 ;
        RECT  6.100 1.860 6.515 2.200 ;
        RECT  1.830 1.060 2.360 2.375 ;
        RECT  2.060 0.595 2.360 2.375 ;
        RECT  1.500 2.375 2.060 2.720 ;
        RECT  6.560 1.055 6.845 1.565 ;
        RECT  6.560 1.335 7.370 1.565 ;
        RECT  10.070 1.915 10.410 2.370 ;
        RECT  9.650 2.140 10.410 2.370 ;
        RECT  7.085 1.335 7.370 3.180 ;
        RECT  9.650 2.140 9.990 3.180 ;
        RECT  7.085 2.950 9.990 3.180 ;
        RECT  10.295 1.095 10.640 1.685 ;
        RECT  9.285 1.455 11.090 1.685 ;
        RECT  9.285 1.455 9.625 1.910 ;
        RECT  10.640 1.455 11.090 1.960 ;
        RECT  10.640 1.455 10.925 2.730 ;
        RECT  9.405 0.635 12.545 0.865 ;
        RECT  9.405 0.635 9.745 1.225 ;
        RECT  8.080 0.995 9.745 1.225 ;
        RECT  8.080 0.995 8.685 1.370 ;
        RECT  12.260 0.635 12.545 2.200 ;
        RECT  8.080 0.995 8.310 2.720 ;
        RECT  7.805 2.380 9.405 2.720 ;
    END
END DFFS_X1_18_SVT_WB

MACRO DFFS_PX8_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFS_PX8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.182  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.455 1.770 0.740 2.200 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.208  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.110 1.695 3.340 2.205 ;
        RECT  2.900 1.695 3.340 2.155 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.195 1.735 13.540 3.175 ;
        RECT  13.200 1.095 13.540 3.175 ;
        RECT  11.880 1.735 13.540 2.100 ;
        RECT  11.880 1.100 12.220 3.175 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.080 0.470 16.420 3.450 ;
        RECT  14.655 1.790 16.420 2.110 ;
        RECT  14.655 0.470 15.180 3.450 ;
        END
    END QN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.227  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.540 1.600 8.910 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.360 4.100 ;
        RECT  16.800 2.475 17.140 4.100 ;
        RECT  15.410 2.640 15.700 4.100 ;
        RECT  13.920 2.695 14.260 4.100 ;
        RECT  11.160 2.695 11.500 4.100 ;
        RECT  8.795 3.515 9.965 4.100 ;
        RECT  4.280 3.515 6.340 4.100 ;
        RECT  2.060 3.515 2.400 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.360 0.180 ;
        RECT  16.800 -0.180 17.140 1.225 ;
        RECT  15.410 -0.180 15.700 1.280 ;
        RECT  11.065 -0.180 11.405 0.405 ;
        RECT  9.460 -0.180 9.800 0.405 ;
        RECT  4.350 -0.180 4.690 0.350 ;
        RECT  2.060 -0.180 2.400 0.350 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.250 1.040 3.800 1.380 ;
        RECT  4.870 1.995 5.210 2.335 ;
        RECT  3.570 2.105 5.210 2.335 ;
        RECT  3.570 1.040 3.800 2.825 ;
        RECT  3.250 2.515 3.800 2.825 ;
        RECT  4.200 1.040 5.825 1.380 ;
        RECT  4.200 1.040 4.540 1.875 ;
        RECT  5.485 1.040 5.825 2.825 ;
        RECT  5.485 2.435 6.705 2.825 ;
        RECT  5.040 2.565 6.705 2.825 ;
        RECT  0.180 1.045 1.270 1.385 ;
        RECT  1.040 1.615 1.600 1.940 ;
        RECT  0.180 2.430 1.270 2.720 ;
        RECT  1.040 1.045 1.270 3.285 ;
        RECT  0.930 2.430 1.270 3.285 ;
        RECT  0.930 3.055 6.910 3.285 ;
        RECT  3.530 3.055 3.870 3.510 ;
        RECT  6.570 3.055 6.910 3.510 ;
        RECT  3.530 0.410 3.870 0.810 ;
        RECT  2.060 0.580 7.850 0.810 ;
        RECT  1.500 1.045 2.360 1.385 ;
        RECT  6.055 0.580 6.285 2.200 ;
        RECT  7.600 0.580 7.850 1.960 ;
        RECT  6.055 1.860 6.515 2.200 ;
        RECT  1.830 1.045 2.360 2.335 ;
        RECT  2.060 0.580 2.360 2.335 ;
        RECT  1.500 2.335 2.060 2.720 ;
        RECT  6.515 1.040 6.800 1.550 ;
        RECT  6.515 1.320 7.370 1.550 ;
        RECT  7.140 1.320 7.370 3.180 ;
        RECT  9.980 1.860 10.265 3.180 ;
        RECT  7.140 2.950 10.265 3.180 ;
        RECT  9.290 1.100 10.780 1.440 ;
        RECT  9.290 1.100 9.630 1.960 ;
        RECT  10.495 1.860 11.650 2.200 ;
        RECT  10.495 1.100 10.780 3.215 ;
        RECT  8.080 0.635 14.425 0.865 ;
        RECT  8.080 0.635 8.430 1.190 ;
        RECT  14.140 0.635 14.425 2.200 ;
        RECT  8.080 0.635 8.310 2.720 ;
        RECT  7.805 2.380 9.410 2.720 ;
    END
END DFFS_PX8_18_SVT_WB

MACRO DFFSR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFSR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.260 2.985 1.830 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.398  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.840 2.380 15.180 3.415 ;
        RECT  14.640 0.870 14.925 3.135 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  16.280 2.385 16.660 3.195 ;
        RECT  16.370 0.580 16.660 3.195 ;
        RECT  16.280 0.580 16.660 1.390 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.229  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.420 1.670 12.760 2.340 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.305  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.780 1.700 11.250 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 17.360 4.100 ;
        RECT  15.560 2.385 15.900 4.100 ;
        RECT  13.620 3.545 13.960 4.100 ;
        RECT  10.780 3.545 12.060 4.100 ;
        RECT  7.580 3.545 7.920 4.100 ;
        RECT  5.560 3.545 5.900 4.100 ;
        RECT  2.240 2.525 2.525 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 17.360 0.180 ;
        RECT  15.615 -0.180 15.900 1.390 ;
        RECT  11.900 -0.180 12.240 0.850 ;
        RECT  6.185 -0.180 6.525 0.815 ;
        RECT  2.400 -0.180 2.740 0.990 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 1.430 1.440 ;
        RECT  1.090 1.100 1.430 2.625 ;
        RECT  0.180 2.395 1.430 2.625 ;
        RECT  0.180 2.395 0.520 2.855 ;
        RECT  3.215 0.970 3.445 2.720 ;
        RECT  4.800 2.565 6.460 2.855 ;
        RECT  4.135 0.970 4.475 1.310 ;
        RECT  4.245 1.505 6.860 1.765 ;
        RECT  6.520 1.505 6.860 1.845 ;
        RECT  4.245 0.970 4.475 2.855 ;
        RECT  4.135 2.515 4.475 2.855 ;
        RECT  4.990 1.995 5.330 2.335 ;
        RECT  4.990 2.105 7.980 2.335 ;
        RECT  7.695 0.970 7.980 2.855 ;
        RECT  6.820 2.105 7.980 2.855 ;
        RECT  6.820 2.515 8.625 2.855 ;
        RECT  8.855 1.765 9.170 2.105 ;
        RECT  8.855 1.765 9.085 3.315 ;
        RECT  4.320 3.085 9.085 3.315 ;
        RECT  4.320 3.085 4.660 3.425 ;
        RECT  3.675 0.410 5.045 0.740 ;
        RECT  7.125 0.410 10.090 0.740 ;
        RECT  4.705 0.410 5.045 1.275 ;
        RECT  7.125 0.410 7.380 1.275 ;
        RECT  4.705 1.045 7.380 1.275 ;
        RECT  8.210 0.410 8.465 1.830 ;
        RECT  1.700 0.680 2.040 2.295 ;
        RECT  9.860 0.410 10.090 2.100 ;
        RECT  3.675 1.860 4.015 2.200 ;
        RECT  1.700 2.060 2.985 2.295 ;
        RECT  2.755 2.060 2.985 3.290 ;
        RECT  3.675 0.410 3.905 3.290 ;
        RECT  2.755 2.950 3.905 3.290 ;
        RECT  1.700 0.680 1.930 3.335 ;
        RECT  1.500 2.995 1.930 3.335 ;
        RECT  8.695 0.970 8.985 1.310 ;
        RECT  8.695 1.035 9.630 1.310 ;
        RECT  9.400 1.035 9.630 3.315 ;
        RECT  9.315 2.515 9.630 3.315 ;
        RECT  13.450 2.050 13.735 3.315 ;
        RECT  9.315 3.085 13.735 3.315 ;
        RECT  13.370 0.970 13.710 1.720 ;
        RECT  12.990 1.380 14.410 1.720 ;
        RECT  11.750 1.540 12.140 1.880 ;
        RECT  14.060 1.380 14.410 1.965 ;
        RECT  11.910 1.540 12.140 2.855 ;
        RECT  12.990 1.380 13.220 2.855 ;
        RECT  11.910 2.570 13.220 2.855 ;
        RECT  12.470 0.410 15.385 0.640 ;
        RECT  10.320 0.970 10.960 1.310 ;
        RECT  12.470 0.410 12.760 1.310 ;
        RECT  10.320 1.080 12.760 1.310 ;
        RECT  15.155 0.410 15.385 1.960 ;
        RECT  15.155 1.620 16.140 1.960 ;
        RECT  10.320 0.970 10.550 2.855 ;
        RECT  9.980 2.515 11.680 2.855 ;
    END
END DFFSR_X4_18_SVT_WB

MACRO DFFSR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFSR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.260 2.985 1.830 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.160 2.420 15.050 2.685 ;
        RECT  14.685 1.050 15.050 2.685 ;
        RECT  14.200 1.050 15.050 1.280 ;
        RECT  14.160 2.420 14.555 3.295 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.720 2.385 16.100 3.210 ;
        RECT  15.810 0.565 16.100 3.210 ;
        RECT  15.775 0.565 16.100 1.390 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.229  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.420 1.670 12.760 2.340 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.305  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.780 1.700 11.250 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  14.960 3.570 15.305 4.100 ;
        RECT  13.420 3.545 13.760 4.100 ;
        RECT  10.780 3.545 12.060 4.100 ;
        RECT  7.580 3.545 7.920 4.100 ;
        RECT  5.560 3.545 5.900 4.100 ;
        RECT  2.240 2.525 2.525 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  14.955 -0.180 15.305 0.350 ;
        RECT  11.900 -0.180 12.240 0.850 ;
        RECT  6.185 -0.180 6.525 0.815 ;
        RECT  2.400 -0.180 2.740 0.990 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 1.430 1.440 ;
        RECT  1.090 1.100 1.430 2.625 ;
        RECT  0.180 2.395 1.430 2.625 ;
        RECT  0.180 2.395 0.520 2.855 ;
        RECT  3.215 0.970 3.445 2.720 ;
        RECT  4.800 2.565 6.460 2.855 ;
        RECT  4.135 0.970 4.475 1.310 ;
        RECT  4.245 1.505 6.860 1.765 ;
        RECT  6.520 1.505 6.860 1.845 ;
        RECT  4.245 0.970 4.475 2.855 ;
        RECT  4.135 2.515 4.475 2.855 ;
        RECT  4.990 1.995 5.330 2.335 ;
        RECT  4.990 2.105 7.980 2.335 ;
        RECT  7.695 0.970 7.980 2.855 ;
        RECT  6.820 2.105 7.980 2.855 ;
        RECT  6.820 2.515 8.625 2.855 ;
        RECT  8.855 1.765 9.170 2.105 ;
        RECT  8.855 1.765 9.085 3.315 ;
        RECT  4.320 3.085 9.085 3.315 ;
        RECT  4.320 3.085 4.660 3.425 ;
        RECT  3.675 0.410 5.045 0.740 ;
        RECT  7.125 0.410 10.090 0.740 ;
        RECT  4.705 0.410 5.045 1.275 ;
        RECT  7.125 0.410 7.380 1.275 ;
        RECT  4.705 1.045 7.380 1.275 ;
        RECT  8.210 0.410 8.465 1.830 ;
        RECT  1.700 0.680 2.040 2.295 ;
        RECT  9.860 0.410 10.090 2.100 ;
        RECT  3.675 1.860 4.015 2.200 ;
        RECT  1.700 2.060 2.985 2.295 ;
        RECT  2.755 2.060 2.985 3.290 ;
        RECT  3.675 0.410 3.905 3.290 ;
        RECT  2.755 2.950 3.905 3.290 ;
        RECT  1.700 0.680 1.930 3.335 ;
        RECT  1.500 2.995 1.930 3.335 ;
        RECT  8.695 0.970 8.985 1.310 ;
        RECT  8.695 1.035 9.630 1.310 ;
        RECT  9.400 1.035 9.630 3.315 ;
        RECT  9.315 2.515 9.630 3.315 ;
        RECT  13.450 2.050 13.735 3.315 ;
        RECT  9.315 3.085 13.735 3.315 ;
        RECT  13.350 1.025 13.730 1.820 ;
        RECT  12.990 1.380 13.730 1.820 ;
        RECT  12.990 1.590 14.455 1.820 ;
        RECT  11.750 1.540 12.140 1.880 ;
        RECT  14.155 1.590 14.455 1.965 ;
        RECT  11.910 1.540 12.140 2.855 ;
        RECT  12.990 1.380 13.220 2.855 ;
        RECT  11.910 2.570 13.220 2.855 ;
        RECT  12.470 0.565 14.825 0.795 ;
        RECT  14.595 0.580 15.535 0.810 ;
        RECT  10.320 0.970 10.960 1.310 ;
        RECT  12.470 0.565 12.760 1.310 ;
        RECT  10.320 1.080 12.760 1.310 ;
        RECT  15.280 0.580 15.535 1.960 ;
        RECT  10.320 0.970 10.550 2.855 ;
        RECT  9.980 2.515 11.680 2.855 ;
    END
END DFFSR_X2_18_SVT_WB

MACRO DFFSR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFSR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.181  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.260 2.985 1.830 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.160 2.420 15.050 2.685 ;
        RECT  14.685 1.050 15.050 2.685 ;
        RECT  14.200 1.050 15.050 1.280 ;
        RECT  14.160 2.420 14.555 2.745 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.720 2.385 16.100 2.745 ;
        RECT  15.810 1.045 16.100 2.745 ;
        RECT  15.775 1.045 16.100 1.390 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.229  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.420 1.670 12.760 2.340 ;
        END
    END RN
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.305  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.780 1.700 11.250 2.150 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  14.960 3.570 15.305 4.100 ;
        RECT  13.420 3.545 13.760 4.100 ;
        RECT  10.780 3.545 12.060 4.100 ;
        RECT  7.580 3.545 7.920 4.100 ;
        RECT  5.560 3.545 5.900 4.100 ;
        RECT  2.240 2.525 2.525 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  14.955 -0.180 15.305 0.350 ;
        RECT  11.900 -0.180 12.240 0.850 ;
        RECT  6.185 -0.180 6.525 0.815 ;
        RECT  2.400 -0.180 2.740 0.990 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 1.430 1.440 ;
        RECT  1.090 1.100 1.430 2.625 ;
        RECT  0.180 2.395 1.430 2.625 ;
        RECT  0.180 2.395 0.520 2.855 ;
        RECT  3.215 0.970 3.445 2.720 ;
        RECT  4.800 2.565 6.460 2.855 ;
        RECT  4.135 0.970 4.475 1.310 ;
        RECT  4.245 1.505 6.860 1.765 ;
        RECT  6.520 1.505 6.860 1.845 ;
        RECT  4.245 0.970 4.475 2.855 ;
        RECT  4.135 2.515 4.475 2.855 ;
        RECT  4.990 1.995 5.330 2.335 ;
        RECT  4.990 2.105 7.980 2.335 ;
        RECT  7.695 0.970 7.980 2.855 ;
        RECT  6.820 2.105 7.980 2.855 ;
        RECT  6.820 2.515 8.625 2.855 ;
        RECT  8.855 1.765 9.170 2.105 ;
        RECT  8.855 1.765 9.085 3.315 ;
        RECT  4.320 3.085 9.085 3.315 ;
        RECT  4.320 3.085 4.660 3.425 ;
        RECT  3.675 0.410 5.045 0.740 ;
        RECT  7.125 0.410 10.090 0.740 ;
        RECT  4.705 0.410 5.045 1.275 ;
        RECT  7.125 0.410 7.380 1.275 ;
        RECT  4.705 1.045 7.380 1.275 ;
        RECT  8.210 0.410 8.465 1.830 ;
        RECT  1.700 0.680 2.040 2.295 ;
        RECT  9.860 0.410 10.090 2.100 ;
        RECT  3.675 1.860 4.015 2.200 ;
        RECT  1.700 2.060 2.985 2.295 ;
        RECT  2.755 2.060 2.985 3.290 ;
        RECT  3.675 0.410 3.905 3.290 ;
        RECT  2.755 2.950 3.905 3.290 ;
        RECT  1.700 0.680 1.930 3.335 ;
        RECT  1.500 2.995 1.930 3.335 ;
        RECT  8.695 0.970 8.985 1.310 ;
        RECT  8.695 1.035 9.630 1.310 ;
        RECT  9.400 1.035 9.630 3.315 ;
        RECT  9.315 2.515 9.630 3.315 ;
        RECT  13.450 2.050 13.735 3.315 ;
        RECT  9.315 3.085 13.735 3.315 ;
        RECT  13.350 1.025 13.730 1.820 ;
        RECT  12.990 1.380 13.730 1.820 ;
        RECT  12.990 1.590 14.455 1.820 ;
        RECT  11.750 1.540 12.140 1.880 ;
        RECT  14.155 1.590 14.455 1.965 ;
        RECT  11.910 1.540 12.140 2.855 ;
        RECT  12.990 1.380 13.220 2.855 ;
        RECT  11.910 2.570 13.220 2.855 ;
        RECT  12.470 0.565 14.825 0.795 ;
        RECT  14.595 0.580 15.535 0.810 ;
        RECT  10.320 0.970 10.960 1.310 ;
        RECT  12.470 0.565 12.760 1.310 ;
        RECT  10.320 1.080 12.760 1.310 ;
        RECT  15.280 0.580 15.535 1.960 ;
        RECT  10.320 0.970 10.550 2.855 ;
        RECT  9.980 2.515 11.680 2.855 ;
    END
END DFFSR_X1_18_SVT_WB

MACRO DFFSQ_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFSQ_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.575 2.260 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.695 1.820 3.275 2.170 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.560 0.535 12.900 3.390 ;
        RECT  11.240 1.665 12.900 2.000 ;
        RECT  11.240 0.535 11.660 3.385 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.201  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.445 0.570 8.970 0.995 ;
        RECT  8.445 0.570 8.740 1.645 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.000 4.100 ;
        RECT  13.280 2.570 13.620 4.100 ;
        RECT  9.510 3.515 10.790 4.100 ;
        RECT  7.800 3.515 8.140 4.100 ;
        RECT  4.440 3.515 5.720 4.100 ;
        RECT  0.780 3.515 2.290 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.000 0.180 ;
        RECT  13.280 -0.180 13.620 1.285 ;
        RECT  9.420 -0.180 10.820 0.405 ;
        RECT  4.360 -0.180 4.700 0.350 ;
        RECT  2.240 -0.180 2.580 0.350 ;
        RECT  0.780 -0.180 1.120 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.230 1.040 3.735 1.325 ;
        RECT  3.505 2.055 5.150 2.300 ;
        RECT  3.505 1.040 3.735 2.825 ;
        RECT  3.230 2.520 3.735 2.825 ;
        RECT  5.000 1.040 5.835 1.825 ;
        RECT  4.140 1.505 5.835 1.825 ;
        RECT  5.555 0.970 5.835 2.825 ;
        RECT  5.480 1.040 5.835 2.825 ;
        RECT  5.480 2.390 6.650 2.825 ;
        RECT  5.000 2.530 6.650 2.825 ;
        RECT  0.220 0.985 1.145 1.425 ;
        RECT  0.805 1.140 1.610 1.480 ;
        RECT  0.220 2.520 1.145 2.860 ;
        RECT  0.805 0.985 1.145 3.285 ;
        RECT  0.805 3.055 6.910 3.285 ;
        RECT  3.470 3.055 3.810 3.510 ;
        RECT  6.570 3.055 6.910 3.510 ;
        RECT  3.460 0.410 3.835 0.810 ;
        RECT  4.995 0.510 7.625 0.740 ;
        RECT  1.530 0.580 5.170 0.810 ;
        RECT  1.530 0.580 2.340 0.910 ;
        RECT  6.065 0.510 6.295 2.120 ;
        RECT  6.065 1.795 6.480 2.120 ;
        RECT  7.395 0.510 7.625 2.210 ;
        RECT  2.020 0.580 2.340 2.340 ;
        RECT  1.830 2.005 2.060 2.825 ;
        RECT  1.530 2.520 2.060 2.825 ;
        RECT  7.930 0.770 8.215 2.730 ;
        RECT  7.800 2.440 8.215 2.730 ;
        RECT  8.600 2.380 8.940 2.730 ;
        RECT  7.800 2.500 8.940 2.730 ;
        RECT  6.525 0.980 7.110 1.325 ;
        RECT  9.740 1.995 10.080 2.320 ;
        RECT  9.170 2.090 10.080 2.320 ;
        RECT  6.880 0.980 7.110 2.730 ;
        RECT  6.880 2.440 7.395 2.730 ;
        RECT  7.165 2.440 7.395 3.285 ;
        RECT  9.170 2.090 9.510 3.285 ;
        RECT  7.165 2.960 9.510 3.285 ;
        RECT  9.980 0.985 10.320 1.630 ;
        RECT  9.980 1.290 10.790 1.630 ;
        RECT  9.070 1.400 10.790 1.630 ;
        RECT  9.070 1.400 9.410 1.860 ;
        RECT  10.450 1.290 10.790 2.890 ;
        RECT  9.980 2.550 10.790 2.890 ;
    END
END DFFSQ_X8_18_SVT_WB

MACRO DFFSQ_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFSQ_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.575 2.260 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.695 1.820 3.275 2.170 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.240 0.535 11.660 3.385 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.201  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.445 0.570 8.970 0.995 ;
        RECT  8.445 0.570 8.740 1.645 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  9.510 3.515 10.790 4.100 ;
        RECT  7.800 3.515 8.140 4.100 ;
        RECT  4.440 3.515 5.720 4.100 ;
        RECT  0.780 3.515 2.290 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  10.480 -0.180 10.820 0.405 ;
        RECT  9.420 -0.180 9.760 0.405 ;
        RECT  4.360 -0.180 4.700 0.350 ;
        RECT  2.240 -0.180 2.580 0.350 ;
        RECT  0.780 -0.180 1.120 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.230 1.040 3.735 1.325 ;
        RECT  3.505 2.055 5.150 2.300 ;
        RECT  3.505 1.040 3.735 2.825 ;
        RECT  3.230 2.520 3.735 2.825 ;
        RECT  5.000 1.040 5.835 1.825 ;
        RECT  4.140 1.505 5.835 1.825 ;
        RECT  5.555 0.970 5.835 2.825 ;
        RECT  5.480 1.040 5.835 2.825 ;
        RECT  5.480 2.390 6.650 2.825 ;
        RECT  5.000 2.530 6.650 2.825 ;
        RECT  0.220 0.985 1.145 1.425 ;
        RECT  0.805 1.140 1.610 1.480 ;
        RECT  0.220 2.520 1.145 2.860 ;
        RECT  0.805 0.985 1.145 3.285 ;
        RECT  0.805 3.055 6.910 3.285 ;
        RECT  3.470 3.055 3.810 3.510 ;
        RECT  6.570 3.055 6.910 3.510 ;
        RECT  3.460 0.410 3.835 0.810 ;
        RECT  4.995 0.510 7.625 0.740 ;
        RECT  1.530 0.580 5.170 0.810 ;
        RECT  1.530 0.580 2.340 0.910 ;
        RECT  6.065 0.510 6.295 2.120 ;
        RECT  6.065 1.795 6.480 2.120 ;
        RECT  7.395 0.510 7.625 2.210 ;
        RECT  2.020 0.580 2.340 2.340 ;
        RECT  1.830 2.005 2.060 2.825 ;
        RECT  1.530 2.520 2.060 2.825 ;
        RECT  7.930 0.770 8.215 2.730 ;
        RECT  7.800 2.440 8.215 2.730 ;
        RECT  8.600 2.380 8.940 2.730 ;
        RECT  7.800 2.500 8.940 2.730 ;
        RECT  6.525 0.980 7.110 1.325 ;
        RECT  9.740 1.995 10.080 2.320 ;
        RECT  9.170 2.090 10.080 2.320 ;
        RECT  6.880 0.980 7.110 2.730 ;
        RECT  6.880 2.440 7.395 2.730 ;
        RECT  7.165 2.440 7.395 3.285 ;
        RECT  9.170 2.090 9.510 3.285 ;
        RECT  7.165 2.960 9.510 3.285 ;
        RECT  9.980 0.985 10.320 1.630 ;
        RECT  9.980 1.290 10.790 1.630 ;
        RECT  9.070 1.400 10.790 1.630 ;
        RECT  9.070 1.400 9.410 1.860 ;
        RECT  10.450 1.290 10.790 2.890 ;
        RECT  9.980 2.550 10.790 2.890 ;
    END
END DFFSQ_X4_18_SVT_WB

MACRO DFFSQ_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFSQ_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.575 2.260 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.695 1.820 3.275 2.170 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.240 0.535 11.620 3.385 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.201  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.445 0.570 8.970 0.995 ;
        RECT  8.445 0.570 8.740 1.645 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  9.510 3.515 10.790 4.100 ;
        RECT  7.800 3.515 8.140 4.100 ;
        RECT  4.440 3.515 5.720 4.100 ;
        RECT  0.780 3.515 2.290 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  9.420 -0.180 10.820 0.405 ;
        RECT  4.360 -0.180 4.700 0.350 ;
        RECT  2.240 -0.180 2.580 0.350 ;
        RECT  0.780 -0.180 1.120 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.230 1.040 3.735 1.325 ;
        RECT  3.505 2.055 5.150 2.300 ;
        RECT  3.505 1.040 3.735 2.825 ;
        RECT  3.230 2.520 3.735 2.825 ;
        RECT  5.000 1.040 5.835 1.825 ;
        RECT  4.140 1.505 5.835 1.825 ;
        RECT  5.555 0.970 5.835 2.825 ;
        RECT  5.480 1.040 5.835 2.825 ;
        RECT  5.480 2.390 6.650 2.825 ;
        RECT  5.000 2.530 6.650 2.825 ;
        RECT  0.220 0.985 1.145 1.425 ;
        RECT  0.805 1.140 1.610 1.480 ;
        RECT  0.220 2.520 1.145 2.860 ;
        RECT  0.805 0.985 1.145 3.285 ;
        RECT  0.805 3.055 6.910 3.285 ;
        RECT  3.470 3.055 3.810 3.510 ;
        RECT  6.570 3.055 6.910 3.510 ;
        RECT  3.460 0.410 3.835 0.810 ;
        RECT  4.995 0.510 7.625 0.740 ;
        RECT  1.530 0.580 5.170 0.810 ;
        RECT  1.530 0.580 2.340 0.910 ;
        RECT  6.065 0.510 6.295 2.120 ;
        RECT  6.065 1.795 6.480 2.120 ;
        RECT  7.395 0.510 7.625 2.210 ;
        RECT  2.020 0.580 2.340 2.340 ;
        RECT  1.830 2.005 2.060 2.825 ;
        RECT  1.530 2.520 2.060 2.825 ;
        RECT  7.930 0.770 8.215 2.730 ;
        RECT  7.800 2.440 8.215 2.730 ;
        RECT  8.600 2.380 8.940 2.730 ;
        RECT  7.800 2.500 8.940 2.730 ;
        RECT  6.525 0.980 7.110 1.325 ;
        RECT  9.740 1.995 10.080 2.320 ;
        RECT  9.170 2.090 10.080 2.320 ;
        RECT  6.880 0.980 7.110 2.730 ;
        RECT  6.880 2.440 7.395 2.730 ;
        RECT  7.165 2.440 7.395 3.285 ;
        RECT  9.170 2.090 9.510 3.285 ;
        RECT  7.165 2.960 9.510 3.285 ;
        RECT  9.980 0.985 10.320 1.630 ;
        RECT  9.980 1.290 10.790 1.630 ;
        RECT  9.070 1.400 10.790 1.630 ;
        RECT  9.070 1.400 9.410 1.860 ;
        RECT  10.450 1.290 10.790 2.890 ;
        RECT  9.980 2.550 10.790 2.890 ;
    END
END DFFSQ_X2_18_SVT_WB

MACRO DFFSQ_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFSQ_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.202  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.575 2.260 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.203  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.695 1.820 3.275 2.170 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.265 0.535 11.620 3.385 ;
        END
    END Q
    PIN SN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.201  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.445 0.570 8.970 0.995 ;
        RECT  8.445 0.570 8.740 1.645 ;
        END
    END SN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  9.510 3.515 10.790 4.100 ;
        RECT  7.800 3.515 8.140 4.100 ;
        RECT  4.440 3.515 5.720 4.100 ;
        RECT  0.780 3.515 2.290 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  9.420 -0.180 10.820 0.405 ;
        RECT  4.360 -0.180 4.700 0.350 ;
        RECT  2.240 -0.180 2.580 0.350 ;
        RECT  0.780 -0.180 1.120 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.230 1.040 3.735 1.325 ;
        RECT  3.505 2.055 5.150 2.300 ;
        RECT  3.505 1.040 3.735 2.825 ;
        RECT  3.230 2.520 3.735 2.825 ;
        RECT  5.000 1.040 5.835 1.825 ;
        RECT  4.140 1.505 5.835 1.825 ;
        RECT  5.555 0.970 5.835 2.825 ;
        RECT  5.480 1.040 5.835 2.825 ;
        RECT  5.480 2.390 6.650 2.825 ;
        RECT  5.000 2.530 6.650 2.825 ;
        RECT  0.220 0.985 1.145 1.425 ;
        RECT  0.805 1.140 1.610 1.480 ;
        RECT  0.220 2.520 1.145 2.860 ;
        RECT  0.805 0.985 1.145 3.285 ;
        RECT  0.805 3.055 6.910 3.285 ;
        RECT  3.470 3.055 3.810 3.510 ;
        RECT  6.570 3.055 6.910 3.510 ;
        RECT  3.460 0.410 3.835 0.810 ;
        RECT  4.995 0.510 7.625 0.740 ;
        RECT  1.530 0.580 5.170 0.810 ;
        RECT  1.530 0.580 2.340 0.910 ;
        RECT  6.065 0.510 6.295 2.120 ;
        RECT  6.065 1.795 6.480 2.120 ;
        RECT  7.395 0.510 7.625 2.210 ;
        RECT  2.020 0.580 2.340 2.340 ;
        RECT  1.830 2.005 2.060 2.825 ;
        RECT  1.530 2.520 2.060 2.825 ;
        RECT  7.930 0.770 8.215 2.730 ;
        RECT  7.800 2.440 8.215 2.730 ;
        RECT  8.600 2.380 8.940 2.730 ;
        RECT  7.800 2.500 8.940 2.730 ;
        RECT  6.525 0.980 7.110 1.325 ;
        RECT  9.740 1.995 10.080 2.320 ;
        RECT  9.170 2.090 10.080 2.320 ;
        RECT  6.880 0.980 7.110 2.730 ;
        RECT  6.880 2.440 7.395 2.730 ;
        RECT  7.165 2.440 7.395 3.285 ;
        RECT  9.170 2.090 9.510 3.285 ;
        RECT  7.165 2.960 9.510 3.285 ;
        RECT  9.980 0.985 10.320 1.630 ;
        RECT  9.980 1.290 10.790 1.630 ;
        RECT  9.070 1.400 10.790 1.630 ;
        RECT  9.070 1.400 9.410 1.860 ;
        RECT  10.450 1.290 10.790 2.890 ;
        RECT  9.980 2.550 10.790 2.890 ;
    END
END DFFSQ_X1_18_SVT_WB

MACRO DFFR_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFR_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.201  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.760 0.745 2.155 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.895 1.720 3.320 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.280 2.080 11.850 2.420 ;
        RECT  11.280 1.100 11.620 3.330 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.800 0.595 13.300 3.330 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 3.250 9.870 3.510 ;
        RECT  6.200 1.905 6.430 3.510 ;
        RECT  4.010 1.905 6.430 2.135 ;
        RECT  4.010 1.795 4.580 2.135 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 14.000 4.100 ;
        RECT  12.040 3.100 12.380 4.100 ;
        RECT  10.105 3.515 10.805 4.100 ;
        RECT  5.630 3.050 5.970 4.100 ;
        RECT  2.070 2.380 2.410 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 14.000 0.180 ;
        RECT  12.040 -0.180 12.380 0.405 ;
        RECT  2.200 -0.180 2.540 0.410 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.080 1.380 1.415 ;
        RECT  1.090 1.080 1.380 2.725 ;
        RECT  0.180 2.385 1.380 2.725 ;
        RECT  4.020 2.365 5.740 2.705 ;
        RECT  3.230 0.875 5.090 1.215 ;
        RECT  4.785 0.875 5.090 1.675 ;
        RECT  4.785 1.440 6.340 1.675 ;
        RECT  3.550 0.875 3.780 2.840 ;
        RECT  3.220 2.500 3.780 2.840 ;
        RECT  5.320 0.875 6.945 1.210 ;
        RECT  6.660 0.875 6.945 3.020 ;
        RECT  1.500 0.540 1.840 0.880 ;
        RECT  2.770 0.410 7.865 0.645 ;
        RECT  1.500 0.640 3.000 0.880 ;
        RECT  1.610 0.640 2.100 2.150 ;
        RECT  7.635 0.410 7.865 2.550 ;
        RECT  7.635 2.210 7.935 2.550 ;
        RECT  1.610 0.540 1.840 3.385 ;
        RECT  1.500 3.045 1.840 3.385 ;
        RECT  9.140 1.545 10.355 1.885 ;
        RECT  7.175 0.920 7.405 3.020 ;
        RECT  9.140 1.545 9.435 3.020 ;
        RECT  7.175 2.780 9.435 3.020 ;
        RECT  8.625 0.945 10.815 1.285 ;
        RECT  10.585 0.945 10.815 3.015 ;
        RECT  8.625 0.945 8.910 2.030 ;
        RECT  10.585 1.860 11.045 3.015 ;
        RECT  9.775 2.675 11.045 3.015 ;
        RECT  8.095 0.485 11.705 0.715 ;
        RECT  11.365 0.635 12.570 0.870 ;
        RECT  8.095 0.485 8.395 1.005 ;
        RECT  12.285 0.635 12.570 1.960 ;
        RECT  8.165 0.485 8.395 2.550 ;
        RECT  8.165 2.260 8.600 2.550 ;
    END
END DFFR_X4_18_SVT_WB

MACRO DFFR_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFR_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.195  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.895 1.720 3.320 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.860 2.380 11.200 2.720 ;
        RECT  10.970 1.100 11.200 2.720 ;
        RECT  10.780 1.100 11.200 1.590 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.360 0.595 12.740 3.330 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 3.250 9.695 3.510 ;
        RECT  6.200 1.910 6.430 3.510 ;
        RECT  4.010 1.910 6.430 2.140 ;
        RECT  4.010 1.800 4.585 2.140 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  11.600 3.100 11.940 4.100 ;
        RECT  10.015 3.515 10.355 4.100 ;
        RECT  5.685 3.050 5.970 4.100 ;
        RECT  2.085 2.380 2.410 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  11.600 -0.180 11.940 0.405 ;
        RECT  2.200 -0.180 2.540 0.350 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.095 1.395 1.380 ;
        RECT  1.090 1.095 1.395 2.820 ;
        RECT  0.180 2.480 1.395 2.820 ;
        RECT  4.025 2.370 5.685 2.655 ;
        RECT  4.025 2.370 4.365 2.975 ;
        RECT  3.220 0.875 5.020 1.215 ;
        RECT  4.785 0.875 5.020 1.680 ;
        RECT  4.785 1.445 6.430 1.680 ;
        RECT  3.550 0.875 3.780 2.755 ;
        RECT  3.220 2.430 3.780 2.755 ;
        RECT  5.250 0.875 6.890 1.215 ;
        RECT  6.660 0.875 6.890 3.020 ;
        RECT  2.765 0.410 7.810 0.645 ;
        RECT  1.500 0.580 2.990 0.890 ;
        RECT  1.625 0.580 2.105 2.150 ;
        RECT  7.580 0.410 7.810 2.515 ;
        RECT  7.580 2.175 7.830 2.515 ;
        RECT  1.625 0.580 1.855 3.385 ;
        RECT  1.500 3.045 1.855 3.385 ;
        RECT  9.035 1.610 10.090 1.950 ;
        RECT  7.120 0.875 7.350 3.020 ;
        RECT  9.035 1.610 9.315 3.020 ;
        RECT  7.120 2.745 9.315 3.020 ;
        RECT  8.520 0.930 10.550 1.215 ;
        RECT  8.520 0.930 8.805 1.830 ;
        RECT  10.320 1.830 10.740 2.170 ;
        RECT  10.320 0.930 10.550 3.015 ;
        RECT  9.545 2.675 10.550 3.015 ;
        RECT  8.040 0.470 11.370 0.700 ;
        RECT  11.030 0.635 12.130 0.870 ;
        RECT  8.040 0.470 8.290 1.075 ;
        RECT  11.845 0.635 12.130 1.960 ;
        RECT  8.060 0.470 8.290 2.500 ;
        RECT  8.060 2.160 8.495 2.500 ;
    END
END DFFR_X2_18_SVT_WB

MACRO DFFR_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFR_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.180  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.885 1.670 3.310 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.840 2.490 11.620 2.830 ;
        RECT  11.005 2.330 11.620 2.830 ;
        RECT  11.005 1.095 11.235 2.830 ;
        RECT  10.840 1.095 11.235 1.430 ;
        END
    END Q
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.360 1.090 12.740 2.830 ;
        END
    END QN
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.275 3.250 9.680 3.510 ;
        RECT  6.275 1.910 6.505 3.510 ;
        RECT  4.010 1.910 6.505 2.140 ;
        RECT  4.010 1.805 4.570 2.140 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  11.600 3.515 11.940 4.100 ;
        RECT  10.340 3.515 10.680 4.100 ;
        RECT  5.760 3.050 6.045 4.100 ;
        RECT  2.115 2.380 2.400 4.100 ;
        RECT  0.740 3.515 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  11.600 -0.180 11.940 0.405 ;
        RECT  2.200 -0.180 2.540 0.350 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 1.425 1.440 ;
        RECT  1.090 1.100 1.425 2.755 ;
        RECT  0.180 2.415 1.425 2.755 ;
        RECT  4.010 2.370 5.760 2.710 ;
        RECT  3.220 0.875 5.080 1.215 ;
        RECT  4.765 0.875 5.080 1.680 ;
        RECT  4.765 1.445 6.490 1.680 ;
        RECT  3.540 0.875 3.770 2.720 ;
        RECT  3.210 2.380 3.770 2.720 ;
        RECT  5.310 0.875 6.965 1.215 ;
        RECT  6.735 0.875 6.965 3.020 ;
        RECT  2.765 0.410 7.925 0.645 ;
        RECT  1.500 0.580 2.990 0.880 ;
        RECT  1.655 0.580 2.100 2.150 ;
        RECT  7.695 0.410 7.925 2.500 ;
        RECT  7.695 2.160 7.990 2.500 ;
        RECT  1.655 0.580 1.885 3.385 ;
        RECT  1.500 3.045 1.885 3.385 ;
        RECT  9.175 1.445 10.125 1.785 ;
        RECT  7.195 0.875 7.465 3.020 ;
        RECT  9.175 1.445 9.405 3.020 ;
        RECT  7.195 2.730 9.405 3.020 ;
        RECT  8.680 0.875 10.585 1.215 ;
        RECT  8.680 0.875 8.945 1.735 ;
        RECT  10.355 1.915 10.775 2.255 ;
        RECT  10.355 0.875 10.585 2.985 ;
        RECT  9.635 2.645 10.585 2.985 ;
        RECT  8.155 0.410 11.370 0.645 ;
        RECT  11.030 0.635 12.130 0.865 ;
        RECT  8.155 0.410 8.450 1.215 ;
        RECT  11.790 0.635 12.130 1.950 ;
        RECT  8.220 0.410 8.450 2.500 ;
        RECT  8.220 2.160 8.560 2.500 ;
    END
END DFFR_X1_18_SVT_WB

MACRO DFFRQ_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFRQ_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.175 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.900 1.770 3.325 2.250 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.300  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.315 0.485 12.655 3.450 ;
        RECT  10.875 1.760 12.655 2.100 ;
        RECT  10.875 0.535 11.215 3.450 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.200 3.240 9.415 3.510 ;
        RECT  6.200 1.920 6.430 3.510 ;
        RECT  4.060 1.920 6.430 2.150 ;
        RECT  4.060 1.770 4.570 2.150 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 13.440 4.100 ;
        RECT  11.550 2.640 11.890 4.100 ;
        RECT  10.110 3.165 10.450 4.100 ;
        RECT  5.685 3.050 5.970 4.100 ;
        RECT  2.140 2.380 2.470 4.100 ;
        RECT  0.810 3.515 1.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 13.440 0.180 ;
        RECT  11.550 -0.180 11.890 1.345 ;
        RECT  10.110 -0.180 10.450 1.225 ;
        RECT  8.220 -0.180 8.560 0.405 ;
        RECT  2.200 -0.180 2.540 0.405 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.095 1.430 1.435 ;
        RECT  1.090 1.095 1.430 2.750 ;
        RECT  0.180 2.410 1.430 2.750 ;
        RECT  4.015 2.380 5.660 2.665 ;
        RECT  4.015 2.380 4.340 2.985 ;
        RECT  3.280 0.875 5.030 1.215 ;
        RECT  4.790 0.875 5.030 1.690 ;
        RECT  4.790 1.445 6.285 1.690 ;
        RECT  3.555 0.875 3.785 2.985 ;
        RECT  3.280 2.645 3.785 2.985 ;
        RECT  5.260 0.875 6.890 1.215 ;
        RECT  6.660 0.875 6.890 3.010 ;
        RECT  1.500 0.535 1.840 0.875 ;
        RECT  2.770 0.410 7.865 0.645 ;
        RECT  1.500 0.635 3.050 0.875 ;
        RECT  1.680 0.635 2.100 2.150 ;
        RECT  7.635 0.410 7.865 2.495 ;
        RECT  7.635 2.205 7.980 2.495 ;
        RECT  1.680 0.635 1.910 3.385 ;
        RECT  1.570 3.045 1.910 3.385 ;
        RECT  8.770 1.915 9.970 2.200 ;
        RECT  7.120 0.875 7.405 3.010 ;
        RECT  8.770 1.915 9.110 3.010 ;
        RECT  7.120 2.725 9.110 3.010 ;
        RECT  9.390 0.690 9.750 1.685 ;
        RECT  8.095 1.455 10.645 1.685 ;
        RECT  8.095 1.455 8.410 1.855 ;
        RECT  10.330 1.455 10.645 2.935 ;
        RECT  9.390 2.640 10.645 2.935 ;
    END
END DFFRQ_X8_18_SVT_WB

MACRO DFFRQ_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFRQ_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.765 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.670 3.365 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.665 0.540 11.085 3.450 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.230 3.250 9.280 3.510 ;
        RECT  6.230 1.920 6.460 3.510 ;
        RECT  4.060 1.920 6.460 2.150 ;
        RECT  4.060 1.770 4.570 2.150 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  9.945 3.180 10.285 4.100 ;
        RECT  5.715 3.050 6.000 4.100 ;
        RECT  2.140 2.380 2.470 4.100 ;
        RECT  0.810 3.515 1.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  9.905 -0.180 10.245 0.405 ;
        RECT  8.215 -0.180 8.555 0.405 ;
        RECT  2.200 -0.180 2.540 0.405 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 1.430 1.440 ;
        RECT  1.090 1.100 1.430 2.750 ;
        RECT  0.180 2.410 1.430 2.750 ;
        RECT  4.055 2.380 5.700 2.665 ;
        RECT  4.055 2.380 4.380 2.985 ;
        RECT  3.280 0.880 5.030 1.220 ;
        RECT  4.790 0.880 5.030 1.690 ;
        RECT  4.790 1.445 6.440 1.690 ;
        RECT  3.595 0.880 3.825 2.720 ;
        RECT  3.280 2.380 3.825 2.720 ;
        RECT  5.260 0.875 6.920 1.215 ;
        RECT  6.690 0.875 6.920 2.945 ;
        RECT  1.500 0.535 1.840 0.875 ;
        RECT  2.770 0.410 7.865 0.645 ;
        RECT  1.500 0.635 3.050 0.875 ;
        RECT  7.635 0.410 7.865 2.425 ;
        RECT  1.680 0.635 2.100 2.150 ;
        RECT  7.635 2.085 7.975 2.425 ;
        RECT  1.680 0.635 1.910 3.385 ;
        RECT  1.570 3.045 1.910 3.385 ;
        RECT  8.610 1.875 9.760 2.200 ;
        RECT  7.150 0.875 7.405 2.995 ;
        RECT  8.610 1.875 8.950 2.995 ;
        RECT  7.150 2.655 8.950 2.995 ;
        RECT  9.405 0.875 9.745 1.645 ;
        RECT  8.095 1.415 10.430 1.645 ;
        RECT  8.095 1.415 8.405 1.755 ;
        RECT  10.090 1.415 10.430 2.950 ;
        RECT  9.180 2.665 10.430 2.950 ;
    END
END DFFRQ_X4_18_SVT_WB

MACRO DFFRQ_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFRQ_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.186  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.685 3.365 2.165 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.680 0.590 11.060 3.395 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.180 3.250 9.350 3.510 ;
        RECT  6.180 1.910 6.410 3.510 ;
        RECT  4.060 1.910 6.410 2.150 ;
        RECT  4.060 1.770 4.570 2.150 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  9.960 3.180 10.300 4.100 ;
        RECT  5.665 3.050 5.950 4.100 ;
        RECT  2.140 2.380 2.470 4.100 ;
        RECT  0.810 3.515 1.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  9.920 -0.180 10.260 0.405 ;
        RECT  8.230 -0.180 8.570 0.405 ;
        RECT  2.200 -0.180 2.540 0.405 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.040 1.430 1.325 ;
        RECT  1.090 1.040 1.430 2.855 ;
        RECT  0.180 2.560 1.430 2.855 ;
        RECT  4.055 2.380 5.665 2.720 ;
        RECT  3.310 0.880 5.050 1.220 ;
        RECT  4.790 0.880 5.050 1.680 ;
        RECT  4.790 1.445 6.410 1.680 ;
        RECT  3.595 0.880 3.825 2.720 ;
        RECT  3.280 2.395 3.825 2.720 ;
        RECT  5.280 0.875 6.875 1.215 ;
        RECT  6.640 0.875 6.875 2.920 ;
        RECT  2.770 0.410 7.880 0.645 ;
        RECT  1.500 0.535 1.910 0.820 ;
        RECT  1.680 0.635 3.080 0.875 ;
        RECT  7.650 0.410 7.880 2.415 ;
        RECT  1.680 0.635 2.100 2.150 ;
        RECT  7.650 2.075 7.990 2.415 ;
        RECT  1.680 0.535 1.910 3.385 ;
        RECT  1.570 3.045 1.910 3.385 ;
        RECT  8.640 1.845 9.760 2.185 ;
        RECT  7.105 0.875 7.420 3.020 ;
        RECT  8.640 1.845 8.970 3.020 ;
        RECT  7.105 2.680 8.970 3.020 ;
        RECT  9.420 0.875 9.760 1.615 ;
        RECT  8.110 1.385 10.450 1.615 ;
        RECT  8.110 1.385 8.420 1.735 ;
        RECT  10.110 1.385 10.450 2.950 ;
        RECT  9.200 2.665 10.450 2.950 ;
    END
END DFFRQ_X2_18_SVT_WB

MACRO DFFRQ_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFRQ_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.185  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.175 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.920 1.720 3.345 2.200 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.680 0.540 11.060 3.295 ;
        END
    END Q
    PIN RN
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.190  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.195 3.245 9.300 3.510 ;
        RECT  6.195 1.920 6.425 3.510 ;
        RECT  4.060 1.920 6.425 2.150 ;
        RECT  4.060 1.770 4.590 2.150 ;
        END
    END RN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  9.960 3.170 10.300 4.100 ;
        RECT  5.680 3.050 5.965 4.100 ;
        RECT  2.150 2.380 2.490 4.100 ;
        RECT  0.810 3.500 1.150 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  9.920 -0.180 10.260 0.410 ;
        RECT  8.230 -0.180 8.570 0.405 ;
        RECT  2.200 -0.180 2.540 0.405 ;
        RECT  0.740 -0.180 1.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.095 1.430 1.435 ;
        RECT  1.090 1.095 1.430 2.815 ;
        RECT  0.180 2.475 1.430 2.815 ;
        RECT  4.035 2.380 5.680 2.665 ;
        RECT  4.035 2.380 4.360 2.985 ;
        RECT  3.300 0.890 5.050 1.230 ;
        RECT  4.810 0.890 5.050 1.690 ;
        RECT  4.810 1.455 6.425 1.690 ;
        RECT  3.575 0.890 3.805 2.985 ;
        RECT  3.300 2.645 3.805 2.985 ;
        RECT  5.280 0.885 6.905 1.225 ;
        RECT  6.655 0.885 6.905 3.015 ;
        RECT  1.500 0.535 1.910 0.875 ;
        RECT  2.770 0.410 7.830 0.655 ;
        RECT  1.500 0.635 3.070 0.875 ;
        RECT  7.600 0.410 7.830 2.445 ;
        RECT  1.680 0.635 2.100 2.155 ;
        RECT  7.600 2.155 7.940 2.445 ;
        RECT  1.680 0.535 1.910 3.370 ;
        RECT  1.570 3.030 1.910 3.370 ;
        RECT  8.330 2.055 9.760 2.340 ;
        RECT  7.135 0.885 7.370 3.015 ;
        RECT  8.330 2.055 8.670 3.015 ;
        RECT  7.135 2.675 8.670 3.015 ;
        RECT  9.420 0.965 9.760 1.825 ;
        RECT  8.060 1.485 10.450 1.825 ;
        RECT  10.110 1.485 10.450 2.940 ;
        RECT  9.200 2.645 10.450 2.940 ;
    END
END DFFRQ_X1_18_SVT_WB

MACRO DFFQ_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFQ_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.745 2.175 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.865 1.450 3.355 2.140 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.300  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  10.315 0.630 10.660 3.325 ;
        RECT  9.000 1.640 10.660 1.995 ;
        RECT  9.000 0.535 9.390 3.325 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.760 4.100 ;
        RECT  11.040 2.480 11.380 4.100 ;
        RECT  7.175 3.515 8.585 4.100 ;
        RECT  4.550 2.705 4.890 4.100 ;
        RECT  2.110 2.415 2.445 4.100 ;
        RECT  0.745 3.515 1.085 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.760 0.180 ;
        RECT  11.040 -0.180 11.380 1.440 ;
        RECT  8.240 -0.180 8.580 0.405 ;
        RECT  6.980 -0.180 7.320 0.750 ;
        RECT  2.205 -0.180 2.545 0.370 ;
        RECT  0.745 -0.180 1.085 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.185 1.095 0.525 1.540 ;
        RECT  0.185 1.310 1.420 1.540 ;
        RECT  1.095 1.310 1.420 2.750 ;
        RECT  0.185 2.410 1.420 2.750 ;
        RECT  3.235 0.880 4.775 1.220 ;
        RECT  4.545 0.880 4.775 1.740 ;
        RECT  4.545 1.400 4.975 1.740 ;
        RECT  3.585 0.880 3.815 3.020 ;
        RECT  3.255 2.680 3.815 3.020 ;
        RECT  5.005 0.880 5.490 1.170 ;
        RECT  4.165 2.135 5.490 2.475 ;
        RECT  5.205 0.880 5.490 3.020 ;
        RECT  5.185 2.135 5.490 3.020 ;
        RECT  5.185 2.675 5.580 3.020 ;
        RECT  1.505 0.535 1.845 0.875 ;
        RECT  2.775 0.410 6.570 0.650 ;
        RECT  1.505 0.600 3.005 0.875 ;
        RECT  1.650 0.600 1.990 2.185 ;
        RECT  1.650 1.845 2.220 2.185 ;
        RECT  6.270 0.410 6.570 2.500 ;
        RECT  1.650 0.600 1.880 3.390 ;
        RECT  1.505 3.050 1.880 3.390 ;
        RECT  5.720 0.880 6.040 1.210 ;
        RECT  6.850 2.085 7.860 2.425 ;
        RECT  5.810 0.880 6.040 3.020 ;
        RECT  6.850 2.085 7.190 3.020 ;
        RECT  5.810 2.730 7.190 3.020 ;
        RECT  7.740 0.880 8.080 1.830 ;
        RECT  6.800 1.490 8.080 1.830 ;
        RECT  6.800 1.600 8.550 1.830 ;
        RECT  8.210 1.600 8.550 3.015 ;
        RECT  7.740 2.675 8.550 3.015 ;
    END
END DFFQ_X8_18_SVT_WB

MACRO DFFQ_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFQ_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.745 2.175 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.865 1.450 3.355 2.140 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.000 0.535 9.390 3.325 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  7.175 3.515 8.585 4.100 ;
        RECT  4.550 2.705 4.890 4.100 ;
        RECT  2.110 2.415 2.445 4.100 ;
        RECT  0.745 3.515 1.085 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  8.240 -0.180 8.580 0.405 ;
        RECT  6.980 -0.180 7.320 0.750 ;
        RECT  2.205 -0.180 2.545 0.370 ;
        RECT  0.745 -0.180 1.085 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.185 1.095 0.525 1.540 ;
        RECT  0.185 1.310 1.420 1.540 ;
        RECT  1.095 1.310 1.420 2.750 ;
        RECT  0.185 2.410 1.420 2.750 ;
        RECT  3.235 0.880 4.775 1.220 ;
        RECT  4.545 0.880 4.775 1.740 ;
        RECT  4.545 1.400 4.975 1.740 ;
        RECT  3.585 0.880 3.815 3.020 ;
        RECT  3.255 2.680 3.815 3.020 ;
        RECT  5.005 0.880 5.490 1.170 ;
        RECT  4.165 2.135 5.490 2.475 ;
        RECT  5.205 0.880 5.490 3.020 ;
        RECT  5.185 2.135 5.490 3.020 ;
        RECT  5.185 2.675 5.580 3.020 ;
        RECT  1.505 0.535 1.845 0.875 ;
        RECT  2.775 0.410 6.570 0.650 ;
        RECT  1.505 0.600 3.005 0.875 ;
        RECT  1.650 0.600 1.990 2.185 ;
        RECT  1.650 1.845 2.220 2.185 ;
        RECT  6.270 0.410 6.570 2.500 ;
        RECT  1.650 0.600 1.880 3.390 ;
        RECT  1.505 3.050 1.880 3.390 ;
        RECT  5.720 0.880 6.040 1.210 ;
        RECT  6.850 2.085 7.860 2.425 ;
        RECT  5.810 0.880 6.040 3.020 ;
        RECT  6.850 2.085 7.190 3.020 ;
        RECT  5.810 2.730 7.190 3.020 ;
        RECT  7.740 0.880 8.080 1.830 ;
        RECT  6.800 1.490 8.080 1.830 ;
        RECT  6.800 1.600 8.550 1.830 ;
        RECT  8.210 1.600 8.550 3.015 ;
        RECT  7.740 2.675 8.550 3.015 ;
    END
END DFFQ_X4_18_SVT_WB

MACRO DFFQ_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFQ_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.760 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.445 3.360 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.000 0.490 9.380 3.370 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  6.610 3.515 8.360 4.100 ;
        RECT  4.490 2.680 4.830 4.100 ;
        RECT  2.110 2.415 2.450 4.100 ;
        RECT  0.740 3.510 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  7.160 -0.180 8.480 0.410 ;
        RECT  2.200 -0.180 2.540 0.400 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.050 0.520 1.420 ;
        RECT  0.180 1.190 1.420 1.420 ;
        RECT  1.090 1.190 1.420 2.735 ;
        RECT  0.180 2.395 1.420 2.735 ;
        RECT  3.260 0.875 4.875 1.215 ;
        RECT  4.640 0.875 4.875 1.750 ;
        RECT  4.640 1.410 4.980 1.750 ;
        RECT  3.695 0.875 4.035 3.020 ;
        RECT  3.260 2.680 4.035 3.020 ;
        RECT  5.105 0.875 5.550 1.215 ;
        RECT  4.265 2.110 5.550 2.450 ;
        RECT  5.210 0.875 5.550 3.020 ;
        RECT  2.770 0.410 6.570 0.645 ;
        RECT  1.500 0.630 3.030 0.970 ;
        RECT  1.650 0.630 1.990 2.180 ;
        RECT  1.650 1.840 2.230 2.180 ;
        RECT  6.285 0.410 6.570 2.520 ;
        RECT  1.650 0.630 1.880 3.390 ;
        RECT  1.500 3.050 1.880 3.390 ;
        RECT  6.950 2.080 7.855 2.380 ;
        RECT  5.780 0.875 6.055 3.040 ;
        RECT  6.950 2.080 7.290 3.040 ;
        RECT  5.780 2.750 7.290 3.040 ;
        RECT  7.740 0.990 8.080 1.850 ;
        RECT  6.800 1.510 8.080 1.850 ;
        RECT  6.800 1.570 8.770 1.850 ;
        RECT  8.430 1.570 8.770 2.950 ;
        RECT  7.740 2.610 8.770 2.950 ;
    END
END DFFQ_X2_18_SVT_WB

MACRO DFFQ_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFQ_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.740 2.150 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.940 1.445 3.360 2.150 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.000 0.515 9.380 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  6.755 3.470 8.505 4.100 ;
        RECT  4.490 2.680 4.830 4.100 ;
        RECT  2.110 2.400 2.450 4.100 ;
        RECT  0.740 3.510 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  7.065 -0.180 8.380 0.405 ;
        RECT  2.200 -0.180 2.540 0.405 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.075 0.520 1.425 ;
        RECT  0.180 1.195 1.420 1.425 ;
        RECT  1.090 1.195 1.420 2.805 ;
        RECT  0.180 2.465 1.420 2.805 ;
        RECT  3.260 0.875 4.865 1.215 ;
        RECT  4.635 0.875 4.865 1.755 ;
        RECT  4.635 1.415 4.980 1.755 ;
        RECT  3.695 0.875 4.035 2.820 ;
        RECT  3.260 2.480 4.035 2.820 ;
        RECT  5.095 0.875 5.440 1.215 ;
        RECT  4.265 2.110 5.440 2.450 ;
        RECT  5.210 0.875 5.440 3.020 ;
        RECT  5.210 2.680 5.550 3.020 ;
        RECT  2.770 0.410 6.570 0.645 ;
        RECT  1.500 0.635 3.030 0.975 ;
        RECT  1.650 0.635 2.100 2.170 ;
        RECT  6.285 0.410 6.570 2.520 ;
        RECT  1.650 0.635 1.880 3.390 ;
        RECT  1.500 3.050 1.880 3.390 ;
        RECT  5.770 0.875 6.055 1.215 ;
        RECT  7.335 2.130 7.840 2.470 ;
        RECT  5.825 0.875 6.055 3.040 ;
        RECT  7.335 2.130 7.565 3.040 ;
        RECT  5.825 2.750 7.565 3.040 ;
        RECT  7.740 0.875 8.080 1.855 ;
        RECT  6.800 1.515 8.770 1.855 ;
        RECT  8.430 1.515 8.770 3.040 ;
        RECT  7.795 2.700 8.770 3.040 ;
    END
END DFFQ_X1_18_SVT_WB

MACRO DFFQN_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFQN_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.745 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.830 1.705 3.245 2.195 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.150  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.000 0.595 9.380 3.330 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  7.350 3.515 8.520 4.100 ;
        RECT  4.430 2.525 4.770 4.100 ;
        RECT  2.105 2.380 2.390 4.100 ;
        RECT  0.740 3.470 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  8.240 -0.180 8.580 0.410 ;
        RECT  6.980 -0.180 7.320 0.750 ;
        RECT  2.200 -0.180 2.540 0.350 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 0.520 1.540 ;
        RECT  0.180 1.310 1.415 1.540 ;
        RECT  1.090 1.310 1.415 2.750 ;
        RECT  0.180 2.410 1.415 2.750 ;
        RECT  3.240 0.880 4.675 1.220 ;
        RECT  4.445 0.880 4.675 1.820 ;
        RECT  4.445 1.480 4.955 1.820 ;
        RECT  3.475 0.880 3.705 2.765 ;
        RECT  3.200 2.425 3.705 2.765 ;
        RECT  5.030 0.880 5.490 1.220 ;
        RECT  3.935 1.955 4.250 2.295 ;
        RECT  3.935 2.050 5.490 2.295 ;
        RECT  5.185 0.880 5.490 2.925 ;
        RECT  5.150 2.050 5.490 2.925 ;
        RECT  2.785 0.410 6.570 0.650 ;
        RECT  1.500 0.580 3.010 0.895 ;
        RECT  1.645 0.580 2.100 2.150 ;
        RECT  6.265 0.410 6.570 2.620 ;
        RECT  1.645 0.580 1.875 3.390 ;
        RECT  1.500 3.050 1.875 3.390 ;
        RECT  7.335 1.915 7.840 2.150 ;
        RECT  5.750 0.880 6.035 3.260 ;
        RECT  7.335 1.915 7.565 3.260 ;
        RECT  5.750 2.920 7.565 3.260 ;
        RECT  7.740 0.880 8.080 1.685 ;
        RECT  6.830 1.400 8.300 1.685 ;
        RECT  8.070 1.345 8.300 2.720 ;
        RECT  7.795 2.380 8.300 2.720 ;
    END
END DFFQN_X4_18_SVT_WB

MACRO DFFQN_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFQN_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.745 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.830 1.705 3.245 2.195 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.022  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.000 0.595 9.380 3.330 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  7.350 3.515 8.520 4.100 ;
        RECT  4.430 2.525 4.770 4.100 ;
        RECT  2.105 2.380 2.390 4.100 ;
        RECT  0.740 3.470 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  8.240 -0.180 8.580 0.410 ;
        RECT  6.980 -0.180 7.320 0.750 ;
        RECT  2.200 -0.180 2.540 0.350 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 0.520 1.540 ;
        RECT  0.180 1.310 1.415 1.540 ;
        RECT  1.090 1.310 1.415 2.750 ;
        RECT  0.180 2.410 1.415 2.750 ;
        RECT  3.240 0.880 4.675 1.220 ;
        RECT  4.445 0.880 4.675 1.820 ;
        RECT  4.445 1.480 4.955 1.820 ;
        RECT  3.475 0.880 3.705 2.765 ;
        RECT  3.200 2.425 3.705 2.765 ;
        RECT  5.030 0.880 5.490 1.220 ;
        RECT  3.935 1.955 4.250 2.295 ;
        RECT  3.935 2.050 5.490 2.295 ;
        RECT  5.185 0.880 5.490 2.985 ;
        RECT  5.150 2.050 5.490 2.985 ;
        RECT  2.785 0.410 6.570 0.650 ;
        RECT  1.500 0.580 3.010 0.895 ;
        RECT  1.645 0.580 2.100 2.150 ;
        RECT  6.265 0.410 6.570 2.620 ;
        RECT  1.645 0.580 1.875 3.390 ;
        RECT  1.500 3.050 1.875 3.390 ;
        RECT  7.335 1.915 7.840 2.150 ;
        RECT  5.750 0.880 6.035 3.085 ;
        RECT  7.335 1.915 7.565 3.085 ;
        RECT  5.750 2.855 7.565 3.085 ;
        RECT  7.740 0.880 8.080 1.685 ;
        RECT  6.830 1.400 8.300 1.685 ;
        RECT  8.070 1.345 8.300 2.720 ;
        RECT  7.795 2.380 8.300 2.720 ;
    END
END DFFQN_X2_18_SVT_WB

MACRO DFFQN_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN DFFQN_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.194  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.745 2.180 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.200  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.830 1.705 3.245 2.195 ;
        END
    END D
    PIN QN
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.000 0.595 9.380 3.330 ;
        END
    END QN
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  7.350 3.515 8.520 4.100 ;
        RECT  4.430 2.645 4.770 4.100 ;
        RECT  2.105 2.380 2.390 4.100 ;
        RECT  0.740 3.470 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  8.240 -0.180 8.580 0.410 ;
        RECT  6.980 -0.180 7.320 0.750 ;
        RECT  2.200 -0.180 2.540 0.350 ;
        RECT  0.740 -0.180 1.080 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 0.520 1.540 ;
        RECT  0.180 1.310 1.415 1.540 ;
        RECT  1.090 1.310 1.415 2.750 ;
        RECT  0.180 2.410 1.415 2.750 ;
        RECT  3.240 0.880 4.675 1.220 ;
        RECT  4.445 0.880 4.675 1.820 ;
        RECT  4.445 1.480 4.955 1.820 ;
        RECT  3.475 0.880 3.705 2.765 ;
        RECT  3.200 2.425 3.705 2.765 ;
        RECT  5.030 0.880 5.490 1.220 ;
        RECT  3.935 1.955 4.250 2.295 ;
        RECT  3.935 2.050 5.490 2.295 ;
        RECT  5.185 0.880 5.490 3.000 ;
        RECT  5.150 2.050 5.490 3.000 ;
        RECT  2.785 0.410 6.570 0.650 ;
        RECT  1.500 0.580 3.010 0.895 ;
        RECT  1.645 0.580 2.100 2.150 ;
        RECT  6.265 0.410 6.570 2.620 ;
        RECT  1.645 0.580 1.875 3.390 ;
        RECT  1.500 3.050 1.875 3.390 ;
        RECT  7.335 1.915 7.840 2.150 ;
        RECT  5.750 0.880 6.035 3.160 ;
        RECT  7.335 1.915 7.565 3.160 ;
        RECT  5.750 2.850 7.565 3.160 ;
        RECT  7.740 0.880 8.080 1.685 ;
        RECT  6.830 1.400 8.300 1.685 ;
        RECT  8.070 1.345 8.300 2.720 ;
        RECT  7.795 2.380 8.300 2.720 ;
    END
END DFFQN_X1_18_SVT_WB

MACRO CLKXOR2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKXOR2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.950 1.915 3.410 2.200 ;
        RECT  1.755 2.380 3.180 2.710 ;
        RECT  2.950 1.915 3.180 2.710 ;
        RECT  0.535 3.185 1.985 3.510 ;
        RECT  1.755 2.380 1.985 3.510 ;
        RECT  0.535 1.620 0.785 3.510 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.070 1.455 4.410 1.940 ;
        RECT  1.790 1.455 4.410 1.685 ;
        RECT  1.790 1.095 2.125 1.685 ;
        RECT  1.510 1.095 2.125 1.405 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.571  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.030 2.380 7.370 3.190 ;
        RECT  6.855 1.065 7.165 2.720 ;
        RECT  5.590 2.380 7.370 2.720 ;
        RECT  5.590 1.065 7.165 1.405 ;
        RECT  5.590 2.380 5.930 3.190 ;
        RECT  5.590 0.630 5.930 1.405 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.775 2.990 8.140 4.100 ;
        RECT  6.315 3.095 6.650 4.100 ;
        RECT  4.310 3.110 4.650 4.100 ;
        RECT  2.215 3.090 2.500 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  6.310 -0.180 6.650 0.815 ;
        RECT  1.870 -0.180 2.210 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.320 0.470 1.245 0.815 ;
        RECT  1.015 1.915 2.720 2.150 ;
        RECT  1.015 0.470 1.245 2.955 ;
        RECT  2.590 0.470 4.650 0.755 ;
        RECT  3.395 0.985 4.875 1.225 ;
        RECT  4.640 1.635 6.625 1.995 ;
        RECT  4.640 0.985 4.875 2.880 ;
        RECT  3.740 2.540 4.875 2.880 ;
        RECT  3.740 2.540 4.040 3.280 ;
        RECT  2.880 2.940 4.040 3.280 ;
    END
END CLKXOR2_X8_18_SVT_WB

MACRO CLKXOR2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKXOR2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.430 1.915 3.890 2.200 ;
        RECT  2.235 2.380 3.660 2.720 ;
        RECT  3.430 1.915 3.660 2.720 ;
        RECT  0.735 3.185 2.465 3.510 ;
        RECT  2.235 2.380 2.465 3.510 ;
        RECT  0.735 1.525 0.985 3.510 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.350 1.455 4.690 1.980 ;
        RECT  2.340 1.455 4.690 1.685 ;
        RECT  2.340 1.095 2.665 1.685 ;
        RECT  1.990 1.095 2.665 1.405 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.914  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.285 1.100 6.585 2.740 ;
        RECT  6.010 0.630 6.350 1.440 ;
        RECT  6.010 2.330 6.335 3.300 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.760 3.160 7.100 4.100 ;
        RECT  5.290 3.160 5.630 4.100 ;
        RECT  4.590 3.110 4.930 4.100 ;
        RECT  2.695 3.090 2.980 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  5.290 -0.180 5.630 0.755 ;
        RECT  2.350 -0.180 2.690 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.520 0.470 0.860 1.165 ;
        RECT  0.520 0.935 1.670 1.165 ;
        RECT  1.405 0.935 1.670 2.150 ;
        RECT  1.405 1.915 3.200 2.150 ;
        RECT  1.405 0.935 1.635 2.955 ;
        RECT  3.070 0.470 4.930 0.755 ;
        RECT  3.790 0.985 5.260 1.225 ;
        RECT  4.920 1.760 6.055 2.100 ;
        RECT  4.920 0.985 5.260 2.880 ;
        RECT  3.995 2.540 5.260 2.880 ;
        RECT  3.995 2.540 4.310 3.450 ;
        RECT  3.360 3.110 4.310 3.450 ;
    END
END CLKXOR2_X4_18_SVT_WB

MACRO CLKXOR2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKXOR2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.480 1.630 3.990 1.970 ;
        RECT  3.480 1.280 3.710 1.970 ;
        RECT  2.950 1.280 3.710 1.510 ;
        RECT  2.950 0.410 3.180 1.510 ;
        RECT  0.700 0.410 3.180 0.640 ;
        RECT  0.700 0.410 0.980 1.730 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 2.200 4.690 2.430 ;
        RECT  4.350 1.860 4.690 2.430 ;
        RECT  1.720 1.760 2.180 2.430 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.848  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.870 2.660 5.460 2.890 ;
        RECT  5.120 1.035 5.460 2.890 ;
        RECT  4.000 1.035 5.460 1.375 ;
        RECT  4.000 0.470 4.340 1.375 ;
        RECT  3.410 0.470 4.340 0.810 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  2.430 2.685 2.770 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.590 -0.180 4.930 0.805 ;
        RECT  0.185 -0.180 0.470 1.210 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.210 0.870 2.720 1.165 ;
        RECT  2.490 0.870 2.720 1.970 ;
        RECT  2.490 1.740 3.250 1.970 ;
        RECT  1.210 0.870 1.440 2.200 ;
        RECT  0.600 1.970 1.440 2.200 ;
        RECT  0.600 1.970 0.940 3.385 ;
        RECT  3.150 3.120 4.930 3.450 ;
    END
END CLKXOR2_X2_18_SVT_WB

MACRO CLKXOR2_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKXOR2_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 1.915 3.320 2.200 ;
        RECT  1.665 2.380 3.090 2.710 ;
        RECT  2.860 1.915 3.090 2.710 ;
        RECT  0.535 2.960 1.895 3.190 ;
        RECT  1.665 2.380 1.895 3.190 ;
        RECT  0.535 1.620 0.785 3.190 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.980 1.455 4.320 1.940 ;
        RECT  1.800 1.455 4.320 1.685 ;
        RECT  1.800 1.095 2.160 1.685 ;
        RECT  1.475 1.095 2.160 1.445 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.352  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.980 2.150 14.320 3.395 ;
        RECT  12.430 1.075 14.320 1.310 ;
        RECT  13.980 0.525 14.320 1.310 ;
        RECT  12.480 2.150 14.320 2.400 ;
        RECT  12.480 2.150 12.820 3.395 ;
        RECT  11.150 0.985 12.820 1.215 ;
        RECT  12.480 0.525 12.820 1.310 ;
        RECT  12.430 0.985 12.775 2.380 ;
        RECT  11.040 2.150 14.320 2.380 ;
        RECT  11.040 2.150 11.380 3.450 ;
        RECT  11.150 0.465 11.380 1.215 ;
        RECT  11.095 0.465 11.380 0.810 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.120 4.100 ;
        RECT  13.200 2.680 13.600 4.100 ;
        RECT  11.760 2.610 12.100 4.100 ;
        RECT  8.945 3.565 9.310 4.100 ;
        RECT  7.685 2.990 8.050 4.100 ;
        RECT  6.225 3.095 6.560 4.100 ;
        RECT  4.220 3.110 4.560 4.100 ;
        RECT  2.125 3.090 2.410 4.100 ;
        RECT  0.180 3.570 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.120 0.180 ;
        RECT  13.240 -0.180 13.595 0.755 ;
        RECT  11.760 -0.180 12.100 0.755 ;
        RECT  8.960 -0.180 9.300 0.350 ;
        RECT  6.410 -0.180 6.750 0.815 ;
        RECT  4.970 -0.180 5.310 0.755 ;
        RECT  1.780 -0.180 2.120 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.320 0.470 1.245 0.815 ;
        RECT  1.015 1.915 2.630 2.150 ;
        RECT  1.015 0.470 1.245 2.730 ;
        RECT  2.500 0.470 4.560 0.755 ;
        RECT  3.305 0.985 4.785 1.225 ;
        RECT  4.550 1.635 6.535 1.995 ;
        RECT  4.550 0.985 4.785 2.880 ;
        RECT  3.650 2.540 4.785 2.880 ;
        RECT  3.650 2.540 3.950 3.280 ;
        RECT  2.790 2.940 3.950 3.280 ;
        RECT  5.690 0.630 6.030 1.405 ;
        RECT  5.690 1.065 7.075 1.405 ;
        RECT  6.765 1.275 9.245 1.585 ;
        RECT  6.765 1.065 7.075 2.720 ;
        RECT  5.500 2.380 7.280 2.720 ;
        RECT  5.500 2.380 5.840 3.190 ;
        RECT  6.940 2.380 7.280 3.190 ;
        RECT  8.175 0.510 8.570 0.810 ;
        RECT  9.715 0.515 10.060 0.810 ;
        RECT  8.175 0.580 10.060 0.810 ;
        RECT  9.720 1.445 11.945 1.685 ;
        RECT  8.400 2.575 10.060 2.805 ;
        RECT  8.400 2.575 8.740 2.880 ;
        RECT  9.720 0.515 10.060 3.395 ;
    END
END CLKXOR2_X16_18_SVT_WB

MACRO CLKXOR2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKXOR2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.240 1.915 3.700 2.200 ;
        RECT  2.045 2.380 3.470 2.720 ;
        RECT  3.240 1.915 3.470 2.720 ;
        RECT  0.735 3.185 2.275 3.510 ;
        RECT  2.045 2.380 2.275 3.510 ;
        RECT  0.735 1.525 0.985 3.510 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.565  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.160 1.455 4.500 1.980 ;
        RECT  2.345 1.455 4.500 1.685 ;
        RECT  2.345 1.095 2.670 1.685 ;
        RECT  1.800 1.095 2.670 1.405 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.604  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.855 2.420 12.185 3.470 ;
        RECT  8.900 2.430 12.185 2.740 ;
        RECT  10.725 2.420 12.185 2.740 ;
        RECT  10.725 0.985 11.095 2.740 ;
        RECT  8.900 0.985 11.095 1.215 ;
        RECT  10.340 2.430 10.680 3.175 ;
        RECT  10.340 0.525 10.680 1.215 ;
        RECT  8.900 2.430 9.240 3.395 ;
        RECT  8.900 0.525 9.240 1.215 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.060 3.150 11.420 4.100 ;
        RECT  9.620 3.115 9.960 4.100 ;
        RECT  8.140 2.635 8.520 4.100 ;
        RECT  6.570 3.160 6.910 4.100 ;
        RECT  5.100 3.160 5.440 4.100 ;
        RECT  4.400 3.110 4.740 4.100 ;
        RECT  2.505 3.090 2.790 4.100 ;
        RECT  0.195 2.515 0.505 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.060 -0.180 11.400 0.755 ;
        RECT  9.620 -0.180 9.960 0.755 ;
        RECT  8.110 -0.180 8.460 0.820 ;
        RECT  5.100 -0.180 5.440 0.755 ;
        RECT  2.160 -0.180 2.500 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.520 0.470 0.860 1.165 ;
        RECT  0.520 0.935 1.480 1.165 ;
        RECT  1.215 0.935 1.480 2.150 ;
        RECT  1.215 1.915 3.010 2.150 ;
        RECT  1.215 0.935 1.445 2.955 ;
        RECT  2.880 0.470 4.740 0.755 ;
        RECT  3.600 0.985 5.070 1.225 ;
        RECT  4.730 1.760 5.865 2.100 ;
        RECT  4.730 0.985 5.070 2.880 ;
        RECT  3.805 2.540 5.070 2.880 ;
        RECT  3.805 2.540 4.120 3.450 ;
        RECT  3.170 3.110 4.120 3.450 ;
        RECT  5.820 0.630 6.160 1.440 ;
        RECT  6.095 1.460 7.160 1.715 ;
        RECT  6.095 1.100 6.395 2.740 ;
        RECT  5.820 2.330 6.145 3.300 ;
        RECT  7.390 1.485 10.410 1.770 ;
        RECT  7.390 0.590 7.730 3.395 ;
    END
END CLKXOR2_X12_18_SVT_WB

MACRO CLKNAND2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKNAND2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.152  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.350 1.820 4.440 2.160 ;
        RECT  1.660 2.135 3.690 2.365 ;
        RECT  1.660 1.860 2.000 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.152  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.280 1.360 5.585 1.960 ;
        RECT  0.870 1.360 5.585 1.590 ;
        RECT  2.660 1.360 3.000 1.905 ;
        RECT  0.870 1.360 3.000 1.630 ;
        RECT  0.520 1.805 1.100 2.145 ;
        RECT  0.870 1.360 1.100 2.145 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.970  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.595 6.045 2.825 ;
        RECT  5.815 0.640 6.045 2.825 ;
        RECT  1.460 0.640 6.045 0.980 ;
        RECT  5.045 2.595 5.400 3.405 ;
        RECT  4.310 0.480 4.685 0.980 ;
        RECT  3.620 2.595 3.960 3.405 ;
        RECT  2.180 2.595 3.960 2.835 ;
        RECT  2.180 2.595 2.520 3.405 ;
        RECT  1.460 0.470 1.815 0.980 ;
        RECT  0.740 2.595 1.075 3.445 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.340 3.065 4.680 4.100 ;
        RECT  2.900 3.065 3.240 4.100 ;
        RECT  1.460 3.065 1.800 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  5.640 -0.180 5.980 0.410 ;
        RECT  2.860 -0.180 3.200 0.390 ;
        RECT  0.180 -0.180 0.520 0.790 ;
        END
    END VSS
END CLKNAND2_X8_18_SVT_WB

MACRO CLKNAND2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKNAND2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.578  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 1.635 2.150 2.140 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.578  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.550 2.370 2.785 2.710 ;
        RECT  2.450 1.860 2.785 2.710 ;
        RECT  0.550 1.860 0.890 2.710 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.524  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.740 2.940 3.245 3.330 ;
        RECT  3.015 1.065 3.245 3.330 ;
        RECT  1.540 1.065 3.245 1.405 ;
        RECT  1.540 0.495 1.880 1.405 ;
        RECT  0.740 2.940 1.080 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.500 3.560 1.840 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.690 -0.180 3.030 0.810 ;
        RECT  0.310 -0.180 0.650 0.810 ;
        END
    END VSS
END CLKNAND2_X4_18_SVT_WB

MACRO CLKNAND2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKNAND2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.175 1.595 1.540 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.510 2.335 1.030 2.675 ;
        RECT  0.510 1.840 0.850 2.675 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.862  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.940 2.905 2.100 3.245 ;
        RECT  1.770 0.470 2.100 3.245 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.700 3.475 2.040 4.100 ;
        RECT  0.220 3.125 0.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.270 -0.180 0.610 0.865 ;
        END
    END VSS
END CLKNAND2_X2_18_SVT_WB

MACRO CLKNAND2_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKNAND2_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.310 2.215 9.045 2.465 ;
        RECT  8.205 1.710 9.045 2.465 ;
        RECT  5.320 1.710 6.145 2.465 ;
        RECT  2.370 1.710 3.280 2.465 ;
        RECT  0.310 1.670 0.875 2.465 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.297  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.565 1.250 9.910 1.600 ;
        RECT  1.260 1.250 9.910 1.480 ;
        RECT  6.520 1.250 7.365 1.590 ;
        RECT  3.870 1.250 4.700 1.605 ;
        RECT  1.260 1.250 1.600 1.600 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.770 2.695 10.500 2.925 ;
        RECT  10.185 0.680 10.500 2.925 ;
        RECT  1.370 0.680 10.500 1.020 ;
        RECT  9.170 2.695 9.510 3.395 ;
        RECT  7.730 2.695 8.070 3.395 ;
        RECT  6.290 2.695 6.630 3.395 ;
        RECT  4.850 2.695 5.190 3.395 ;
        RECT  3.355 2.695 3.750 3.395 ;
        RECT  2.080 2.695 2.485 3.395 ;
        RECT  0.770 2.695 1.145 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.640 4.100 ;
        RECT  8.450 3.180 8.790 4.100 ;
        RECT  7.010 3.180 7.350 4.100 ;
        RECT  5.570 3.180 5.910 4.100 ;
        RECT  4.130 3.180 4.470 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.640 0.180 ;
        RECT  8.610 -0.180 8.950 0.410 ;
        RECT  2.560 -0.180 2.900 0.450 ;
        END
    END VSS
END CLKNAND2_X16_18_SVT_WB

MACRO CLKNAND2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKNAND2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.725  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.460 2.135 6.080 2.365 ;
        RECT  5.690 1.555 6.080 2.365 ;
        RECT  2.860 1.555 3.200 2.365 ;
        RECT  0.460 1.860 0.800 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.725  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.920 1.095 7.260 1.835 ;
        RECT  1.900 1.095 7.260 1.325 ;
        RECT  4.060 1.095 4.400 1.795 ;
        RECT  1.900 1.095 2.240 1.795 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.940 2.640 7.725 2.870 ;
        RECT  7.490 0.635 7.725 2.870 ;
        RECT  0.220 0.635 7.725 0.865 ;
        RECT  6.700 2.640 7.040 3.450 ;
        RECT  0.940 2.640 7.040 2.880 ;
        RECT  5.940 0.470 6.365 0.865 ;
        RECT  5.260 2.640 5.600 3.450 ;
        RECT  3.820 2.640 4.160 3.450 ;
        RECT  3.070 0.500 3.480 0.865 ;
        RECT  2.380 2.640 2.720 3.450 ;
        RECT  0.940 2.640 1.280 3.450 ;
        RECT  0.220 0.470 0.580 0.865 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.980 3.110 6.320 4.100 ;
        RECT  4.540 3.110 4.880 4.100 ;
        RECT  3.100 3.110 3.440 4.100 ;
        RECT  1.660 3.110 2.000 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  7.170 -0.180 7.510 0.405 ;
        RECT  4.500 -0.180 4.840 0.405 ;
        RECT  1.700 -0.180 2.040 0.405 ;
        END
    END VSS
END CLKNAND2_X12_18_SVT_WB

MACRO CLKMUX2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKMUX2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.060 1.640 4.530 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.830 1.590 2.660 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.571  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.620 2.570 6.950 3.390 ;
        RECT  6.290 0.585 6.635 2.800 ;
        RECT  5.190 2.570 6.950 2.800 ;
        RECT  5.190 0.585 6.635 0.815 ;
        RECT  5.190 0.475 5.560 0.815 ;
        RECT  5.190 2.570 5.530 3.390 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.472  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.590 1.260 2.875 1.960 ;
        RECT  0.575 1.260 2.875 1.600 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.910 3.110 6.265 4.100 ;
        RECT  4.430 2.440 4.770 4.100 ;
        RECT  0.960 3.515 1.300 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.950 -0.180 6.290 0.350 ;
        RECT  4.430 -0.180 4.770 0.755 ;
        RECT  1.000 -0.180 1.340 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.470 0.620 0.810 ;
        RECT  0.115 0.470 0.345 3.230 ;
        RECT  1.910 1.860 2.195 3.230 ;
        RECT  0.115 2.890 2.195 3.230 ;
        RECT  3.575 1.860 3.830 3.230 ;
        RECT  0.115 3.000 3.830 3.230 ;
        RECT  3.105 1.135 5.225 1.395 ;
        RECT  4.905 1.135 5.225 1.960 ;
        RECT  4.905 1.665 5.855 1.960 ;
        RECT  3.105 0.470 3.345 2.720 ;
        RECT  2.425 2.380 3.345 2.720 ;
    END
END CLKMUX2_X8_18_SVT_WB

MACRO CLKMUX2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKMUX2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.055 1.120 4.485 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.000 1.190 1.555 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.612  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.720 2.235 7.140 3.235 ;
        RECT  6.795 1.010 7.140 3.235 ;
        RECT  5.280 1.010 7.140 1.240 ;
        RECT  5.280 2.235 7.140 2.465 ;
        RECT  5.280 2.235 5.620 3.235 ;
        RECT  5.280 0.505 5.620 1.240 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.690 2.545 3.365 2.775 ;
        RECT  3.045 1.765 3.365 2.775 ;
        RECT  0.690 1.840 1.090 2.775 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.000 2.695 6.340 4.100 ;
        RECT  4.520 3.515 4.860 4.100 ;
        RECT  0.985 3.515 1.325 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  4.520 -0.180 4.860 0.405 ;
        RECT  0.985 -0.180 1.325 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.185 0.635 2.515 0.915 ;
        RECT  0.225 0.575 0.565 0.930 ;
        RECT  2.160 0.635 2.515 1.435 ;
        RECT  2.160 1.095 3.825 1.435 ;
        RECT  2.160 0.635 2.510 2.120 ;
        RECT  0.185 0.580 0.415 3.295 ;
        RECT  0.185 3.010 0.600 3.295 ;
        RECT  3.290 0.465 3.630 0.865 ;
        RECT  3.290 0.635 5.050 0.865 ;
        RECT  4.715 0.635 5.050 3.285 ;
        RECT  2.625 3.005 5.050 3.285 ;
        RECT  2.625 3.005 3.630 3.345 ;
    END
END CLKMUX2_X6_18_SVT_WB

MACRO CLKMUX2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKMUX2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.730 1.095 4.415 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.860 1.160 1.650 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.135  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.135 0.495 5.530 3.280 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.715 2.175 3.380 2.405 ;
        RECT  2.830 1.725 3.380 2.405 ;
        RECT  0.715 1.845 0.945 2.405 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.225 2.630 4.600 4.100 ;
        RECT  0.940 2.970 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.055 -0.180 4.690 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.575 0.520 0.915 ;
        RECT  0.180 0.635 2.275 0.915 ;
        RECT  1.880 0.635 2.275 1.435 ;
        RECT  1.880 1.095 3.345 1.435 ;
        RECT  1.880 0.635 2.265 1.925 ;
        RECT  0.180 0.575 0.485 3.295 ;
        RECT  2.820 0.525 3.160 0.865 ;
        RECT  2.820 0.635 4.905 0.865 ;
        RECT  4.675 0.635 4.905 2.290 ;
        RECT  3.670 2.060 4.905 2.290 ;
        RECT  3.670 2.060 3.900 3.285 ;
        RECT  2.175 3.010 3.900 3.285 ;
    END
END CLKMUX2_X4_18_SVT_WB

MACRO CLKMUX2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKMUX2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.237  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.345 1.750 4.065 2.115 ;
        RECT  3.655 1.095 4.065 2.115 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.237  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.025 1.210 1.720 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.678  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.775 3.010 5.480 3.385 ;
        RECT  5.150 0.480 5.480 3.385 ;
        RECT  4.775 0.480 5.480 0.820 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.388  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.535 2.955 2.765 ;
        RECT  2.595 1.765 2.955 2.765 ;
        RECT  0.650 1.925 1.025 2.765 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.075 3.515 4.415 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.075 -0.180 4.415 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 0.495 0.510 0.915 ;
        RECT  0.140 0.635 2.615 0.915 ;
        RECT  2.315 0.635 2.615 1.435 ;
        RECT  2.315 1.095 3.425 1.435 ;
        RECT  1.950 1.195 3.425 1.435 ;
        RECT  1.950 1.195 2.265 2.125 ;
        RECT  0.140 0.495 0.415 3.295 ;
        RECT  0.140 3.005 0.555 3.295 ;
        RECT  2.845 0.460 3.185 0.865 ;
        RECT  2.845 0.635 4.545 0.865 ;
        RECT  4.295 0.635 4.545 3.285 ;
        RECT  2.325 3.005 4.545 3.285 ;
        RECT  2.325 3.005 3.185 3.345 ;
    END
END CLKMUX2_X3_18_SVT_WB

MACRO CLKMUX2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKMUX2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.930 1.095 4.340 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.060 1.100 1.705 1.540 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.768  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.080 0.470 5.460 3.385 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.445  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.685 2.500 3.185 2.730 ;
        RECT  2.900 1.750 3.185 2.730 ;
        RECT  0.685 1.770 1.035 2.730 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.320 3.515 4.660 4.100 ;
        RECT  0.965 3.515 1.305 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.320 -0.180 4.660 0.405 ;
        RECT  0.965 -0.180 1.305 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.165 0.470 0.545 0.870 ;
        RECT  0.165 0.640 2.860 0.870 ;
        RECT  2.560 0.640 2.860 1.405 ;
        RECT  2.560 1.095 3.680 1.405 ;
        RECT  1.935 1.100 3.680 1.405 ;
        RECT  1.935 1.100 2.225 2.035 ;
        RECT  0.165 0.470 0.400 3.295 ;
        RECT  0.165 2.960 0.545 3.295 ;
        RECT  3.090 0.525 3.430 0.865 ;
        RECT  3.090 0.635 4.850 0.865 ;
        RECT  4.570 0.635 4.850 3.285 ;
        RECT  2.595 3.010 4.850 3.285 ;
        RECT  2.595 3.010 3.430 3.350 ;
    END
END CLKMUX2_X2_18_SVT_WB

MACRO CLKMUX2_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKMUX2_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.895 1.095 3.325 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.625 1.210 1.495 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.328  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.655 1.225 11.695 1.600 ;
        RECT  11.320 0.470 11.695 1.600 ;
        RECT  11.120 1.225 11.460 3.135 ;
        RECT  8.255 0.600 10.270 0.830 ;
        RECT  9.885 0.485 10.270 0.830 ;
        RECT  9.680 0.600 10.020 3.135 ;
        RECT  8.255 2.320 10.020 2.665 ;
        RECT  9.655 0.600 10.020 2.665 ;
        RECT  8.255 0.485 8.590 0.830 ;
        RECT  8.255 2.320 8.580 3.190 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.349  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.685 1.915 2.205 2.150 ;
        RECT  1.775 1.765 2.205 2.150 ;
        RECT  0.685 1.915 1.025 2.255 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  10.400 2.395 10.740 4.100 ;
        RECT  8.960 2.895 9.300 4.100 ;
        RECT  4.840 2.575 5.180 4.100 ;
        RECT  3.360 3.515 3.700 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  10.620 -0.180 10.960 0.770 ;
        RECT  9.000 -0.180 9.340 0.350 ;
        RECT  7.520 -0.180 7.860 0.815 ;
        RECT  6.355 -0.180 6.700 0.350 ;
        RECT  4.840 -0.180 5.180 1.345 ;
        RECT  3.360 -0.180 3.700 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.575 0.520 0.915 ;
        RECT  0.180 0.635 1.955 0.915 ;
        RECT  1.725 0.635 1.955 1.435 ;
        RECT  1.725 1.095 2.665 1.435 ;
        RECT  1.905 2.435 2.665 2.775 ;
        RECT  2.435 1.095 2.665 2.775 ;
        RECT  0.180 2.545 2.665 2.775 ;
        RECT  0.180 2.545 0.520 3.295 ;
        RECT  2.185 0.525 2.470 0.865 ;
        RECT  2.185 0.635 3.785 0.865 ;
        RECT  3.555 0.635 3.785 3.285 ;
        RECT  2.130 3.005 3.785 3.285 ;
        RECT  2.130 3.005 2.470 3.345 ;
        RECT  4.090 1.665 6.265 1.950 ;
        RECT  4.090 0.535 4.460 3.385 ;
        RECT  5.600 0.475 5.940 1.295 ;
        RECT  5.600 0.955 6.860 1.295 ;
        RECT  6.495 1.265 9.280 1.615 ;
        RECT  6.495 0.955 6.860 2.920 ;
        RECT  5.600 2.570 7.260 2.920 ;
        RECT  5.600 2.570 5.940 3.390 ;
        RECT  6.920 2.570 7.260 3.390 ;
    END
END CLKMUX2_X16_18_SVT_WB

MACRO CLKMUX2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKMUX2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.237  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.345 1.750 4.065 2.115 ;
        RECT  3.655 1.095 4.065 2.115 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.237  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.025 1.210 1.720 1.590 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.611  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.795 2.545 12.140 3.310 ;
        RECT  8.880 2.545 12.140 2.785 ;
        RECT  10.445 0.530 10.815 0.860 ;
        RECT  10.360 2.545 10.700 3.390 ;
        RECT  10.185 0.635 10.565 2.785 ;
        RECT  8.920 0.635 10.565 0.865 ;
        RECT  8.880 2.545 9.285 3.350 ;
        RECT  8.920 0.530 9.270 0.865 ;
        END
    END Q
    PIN S0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.388  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.535 2.955 2.765 ;
        RECT  2.595 1.765 2.955 2.765 ;
        RECT  0.650 1.925 1.025 2.765 ;
        END
    END S0
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.080 3.065 11.420 4.100 ;
        RECT  9.640 3.105 9.980 4.100 ;
        RECT  8.255 2.565 8.485 4.100 ;
        RECT  4.075 3.515 4.415 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.185 -0.180 11.545 0.875 ;
        RECT  9.685 -0.180 10.035 0.350 ;
        RECT  8.190 -0.180 8.560 0.775 ;
        RECT  5.645 -0.180 5.985 1.290 ;
        RECT  4.075 -0.180 4.415 0.405 ;
        RECT  0.940 -0.180 1.280 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 0.495 0.510 0.915 ;
        RECT  0.140 0.635 2.615 0.915 ;
        RECT  2.315 0.635 2.615 1.435 ;
        RECT  2.315 1.095 3.425 1.435 ;
        RECT  1.950 1.195 3.425 1.435 ;
        RECT  1.950 1.195 2.265 2.125 ;
        RECT  0.140 0.495 0.415 3.295 ;
        RECT  0.140 3.005 0.555 3.295 ;
        RECT  2.845 0.460 3.185 0.865 ;
        RECT  2.845 0.635 4.545 0.865 ;
        RECT  4.295 0.635 4.545 3.285 ;
        RECT  2.325 3.005 4.545 3.285 ;
        RECT  2.325 3.005 3.185 3.345 ;
        RECT  4.775 0.480 5.320 0.820 ;
        RECT  5.025 1.620 6.820 1.950 ;
        RECT  5.025 0.480 5.320 3.385 ;
        RECT  4.775 3.010 5.320 3.385 ;
        RECT  6.405 0.465 6.745 1.290 ;
        RECT  6.405 1.015 7.360 1.290 ;
        RECT  7.050 1.200 9.955 1.550 ;
        RECT  7.050 1.015 7.360 2.660 ;
        RECT  6.155 2.380 7.815 2.660 ;
        RECT  6.155 2.380 6.495 3.190 ;
        RECT  7.475 2.380 7.815 3.190 ;
    END
END CLKMUX2_X12_18_SVT_WB

MACRO CLKINV_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.048  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.615 1.665 1.565 2.160 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.571  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.570 2.560 3.390 ;
        RECT  0.900 2.570 2.560 2.920 ;
        RECT  1.795 1.000 2.160 2.920 ;
        RECT  0.900 1.000 2.160 1.295 ;
        RECT  0.900 2.570 1.240 3.390 ;
        RECT  0.900 0.475 1.240 1.295 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.180 2.580 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.660 -0.180 2.000 0.765 ;
        RECT  0.180 -0.180 0.520 0.825 ;
        END
    END VSS
END CLKINV_X8_18_SVT_WB

MACRO CLKINV_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.786  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.540 1.620 1.565 2.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.923  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.220 2.380 2.560 3.190 ;
        RECT  0.900 2.380 2.560 2.660 ;
        RECT  1.795 1.015 2.105 2.660 ;
        RECT  0.900 1.015 2.105 1.290 ;
        RECT  0.900 2.380 1.240 3.190 ;
        RECT  0.900 0.465 1.240 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.600 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.180 -0.180 0.520 1.290 ;
        END
    END VSS
END CLKINV_X6_18_SVT_WB

MACRO CLKINV_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.524  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.215 1.440 1.645 2.320 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.914  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.905 2.695 1.245 3.205 ;
        RECT  0.700 0.605 1.245 0.890 ;
        RECT  0.700 0.605 0.985 2.925 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.625 3.110 1.965 4.100 ;
        RECT  0.185 3.110 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.185 -0.180 0.470 0.945 ;
        END
    END VSS
END CLKINV_X4_18_SVT_WB

MACRO CLKINV_X40_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X40_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 5.096  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.155 5.400 1.680 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.817  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.900 0.580 10.315 0.830 ;
        RECT  9.945 0.525 10.315 0.830 ;
        RECT  9.540 1.945 9.880 3.150 ;
        RECT  0.900 1.965 9.880 2.205 ;
        RECT  5.660 1.945 9.880 2.205 ;
        RECT  8.430 0.525 8.795 0.830 ;
        RECT  8.100 1.945 8.440 3.135 ;
        RECT  6.920 0.525 7.260 0.830 ;
        RECT  6.660 1.945 7.000 3.135 ;
        RECT  5.660 0.580 6.030 2.205 ;
        RECT  5.480 0.525 5.820 0.830 ;
        RECT  5.220 1.965 5.560 3.135 ;
        RECT  4.040 0.525 4.380 0.830 ;
        RECT  3.780 1.965 4.120 3.135 ;
        RECT  2.515 0.530 2.860 0.830 ;
        RECT  2.340 1.965 2.680 3.135 ;
        RECT  0.900 1.965 1.240 3.135 ;
        RECT  0.900 0.525 1.240 0.830 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  10.260 2.435 10.600 4.100 ;
        RECT  8.820 2.435 9.160 4.100 ;
        RECT  7.380 2.435 7.720 4.100 ;
        RECT  5.940 2.435 6.280 4.100 ;
        RECT  4.500 2.435 4.840 4.100 ;
        RECT  3.060 2.435 3.400 4.100 ;
        RECT  1.620 2.435 1.960 4.100 ;
        RECT  0.180 2.435 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  10.680 -0.180 11.020 0.765 ;
        RECT  9.200 -0.180 9.540 0.350 ;
        RECT  7.680 -0.180 8.020 0.350 ;
        RECT  3.280 -0.180 3.620 0.350 ;
        RECT  1.700 -0.180 2.050 0.350 ;
        RECT  0.180 -0.180 0.520 0.765 ;
        END
    END VSS
END CLKINV_X40_18_SVT_WB

MACRO CLKINV_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.389  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.215 1.440 1.645 2.320 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.676  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.905 2.695 1.245 3.205 ;
        RECT  0.700 0.525 1.245 0.810 ;
        RECT  0.700 0.525 0.985 2.925 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.625 3.110 1.965 4.100 ;
        RECT  0.185 3.110 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.185 -0.180 0.470 0.865 ;
        END
    END VSS
END CLKINV_X3_18_SVT_WB

MACRO CLKINV_X32_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X32_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 4.193  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.205 4.100 1.650 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.548  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.965 0.580 9.090 0.860 ;
        RECT  8.740 0.475 9.090 0.860 ;
        RECT  0.965 0.580 8.495 0.865 ;
        RECT  8.150 1.940 8.490 3.135 ;
        RECT  0.965 1.940 8.490 2.205 ;
        RECT  7.210 0.535 7.550 0.865 ;
        RECT  6.710 1.940 7.050 3.135 ;
        RECT  5.690 0.535 6.030 0.865 ;
        RECT  5.270 1.940 5.610 3.135 ;
        RECT  4.530 0.580 4.950 2.205 ;
        RECT  4.170 0.535 4.510 0.865 ;
        RECT  3.830 1.940 4.170 3.135 ;
        RECT  2.650 0.535 2.990 0.865 ;
        RECT  2.390 1.940 2.730 3.135 ;
        RECT  0.965 1.940 1.290 3.200 ;
        RECT  0.965 0.480 1.290 0.865 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  8.870 2.435 9.210 4.100 ;
        RECT  7.430 2.435 7.770 4.100 ;
        RECT  5.990 2.435 6.330 4.100 ;
        RECT  4.550 2.435 4.890 4.100 ;
        RECT  3.110 2.435 3.450 4.100 ;
        RECT  1.670 2.435 2.010 4.100 ;
        RECT  0.230 2.435 0.570 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  7.985 -0.180 8.325 0.350 ;
        RECT  6.450 -0.180 6.790 0.350 ;
        RECT  4.930 -0.180 5.270 0.350 ;
        RECT  3.410 -0.180 3.750 0.350 ;
        RECT  1.750 -0.180 2.100 0.350 ;
        RECT  0.230 -0.180 0.570 0.785 ;
        END
    END VSS
END CLKINV_X32_18_SVT_WB

MACRO CLKINV_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.341  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.210 0.985 1.995 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.590 1.540 3.295 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  0.440 2.400 0.780 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  0.180 -0.180 0.520 0.980 ;
        END
    END VSS
END CLKINV_X2_18_SVT_WB

MACRO CLKINV_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 3.149  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.115 3.570 1.665 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.049  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.675 1.975 7.015 3.135 ;
        RECT  0.915 1.975 7.015 2.205 ;
        RECT  0.915 0.585 5.955 0.815 ;
        RECT  5.615 0.555 5.955 0.815 ;
        RECT  5.235 1.975 5.575 3.135 ;
        RECT  4.095 0.555 4.435 0.815 ;
        RECT  4.035 0.585 4.370 2.205 ;
        RECT  3.795 1.975 4.135 3.135 ;
        RECT  2.575 0.555 2.915 0.815 ;
        RECT  2.355 1.975 2.695 3.135 ;
        RECT  0.915 1.975 1.255 3.145 ;
        RECT  0.915 0.530 1.255 0.815 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.955 2.435 6.295 4.100 ;
        RECT  4.515 2.435 4.855 4.100 ;
        RECT  3.075 2.435 3.415 4.100 ;
        RECT  1.635 2.435 1.975 4.100 ;
        RECT  0.195 2.435 0.535 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.335 -0.180 6.675 0.785 ;
        RECT  4.855 -0.180 5.195 0.355 ;
        RECT  3.335 -0.180 3.675 0.355 ;
        RECT  1.815 -0.180 2.155 0.355 ;
        RECT  0.180 -0.180 0.520 0.785 ;
        END
    END VSS
END CLKINV_X24_18_SVT_WB

MACRO CLKINV_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.620  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.155 0.685 1.675 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.100  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.980 0.495 5.320 3.150 ;
        RECT  0.915 1.135 5.320 1.595 ;
        RECT  3.540 0.540 3.880 3.135 ;
        RECT  2.220 0.540 2.560 3.135 ;
        RECT  0.915 0.485 1.240 3.190 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  4.260 2.375 4.600 4.100 ;
        RECT  0.180 2.435 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.260 -0.180 4.600 0.820 ;
        RECT  0.180 -0.180 0.520 0.775 ;
        END
    END VSS
END CLKINV_X20_18_SVT_WB

MACRO CLKINV_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.347  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.605 1.210 0.985 1.745 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.634  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.215 0.590 1.540 3.075 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.680 4.100 ;
        RECT  0.440 2.890 0.780 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.680 0.180 ;
        RECT  0.180 -0.180 0.520 0.980 ;
        END
    END VSS
END CLKINV_X1_18_SVT_WB

MACRO CLKINV_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.037  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.125 0.735 1.660 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.328  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.830 0.540 4.170 3.135 ;
        RECT  0.965 1.225 4.170 1.600 ;
        RECT  2.390 0.495 2.730 3.135 ;
        RECT  0.965 1.220 2.730 1.600 ;
        RECT  0.965 0.485 1.290 3.190 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.110 2.395 3.450 4.100 ;
        RECT  1.670 2.395 2.010 4.100 ;
        RECT  0.230 2.395 0.570 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.110 -0.180 3.450 0.770 ;
        RECT  1.670 -0.180 2.010 0.775 ;
        RECT  0.230 -0.180 0.570 0.815 ;
        END
    END VSS
END CLKINV_X16_18_SVT_WB

MACRO CLKINV_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKINV_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.567  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.200 2.040 1.790 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.611  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.860 2.545 4.120 2.785 ;
        RECT  2.365 0.590 2.785 2.785 ;
        RECT  2.405 0.530 2.785 2.785 ;
        RECT  2.340 2.545 2.680 3.390 ;
        RECT  0.900 0.590 2.785 0.865 ;
        RECT  0.900 0.530 1.260 0.865 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.060 3.065 3.400 4.100 ;
        RECT  1.620 3.105 1.960 4.100 ;
        RECT  0.235 2.565 0.465 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.165 -0.180 3.525 0.875 ;
        RECT  1.650 -0.180 2.025 0.350 ;
        RECT  0.170 -0.180 0.540 0.775 ;
        END
    END VSS
END CLKINV_X12_18_SVT_WB

MACRO CLKBUF_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.436  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.675 0.840 2.170 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.877  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 0.700 3.885 3.395 ;
        RECT  3.560 0.460 3.885 3.395 ;
        RECT  2.060 2.225 3.885 2.465 ;
        RECT  2.060 0.700 3.885 0.935 ;
        RECT  2.060 2.225 2.400 3.395 ;
        RECT  2.060 0.490 2.400 0.935 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  2.780 2.695 3.120 4.100 ;
        RECT  0.170 3.560 0.530 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  2.820 -0.180 3.160 0.470 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.715 1.065 1.330 1.400 ;
        RECT  0.715 0.460 1.085 1.400 ;
        RECT  1.070 1.295 3.270 1.590 ;
        RECT  1.070 1.295 1.345 2.915 ;
        RECT  0.740 2.575 1.345 2.915 ;
    END
END CLKBUF_X8_18_SVT_WB

MACRO CLKBUF_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.210 0.625 2.165 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.070  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.535 1.920 2.125 2.855 ;
        RECT  1.635 0.505 2.125 2.855 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.955 3.565 1.295 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.355 -0.180 2.695 0.795 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 0.475 1.405 0.830 ;
        RECT  1.075 0.475 1.405 1.520 ;
        RECT  1.075 0.475 1.305 2.815 ;
        RECT  0.165 2.490 1.305 2.815 ;
        RECT  0.165 2.490 0.545 3.330 ;
    END
END CLKBUF_X6_18_SVT_WB

MACRO CLKBUF_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.358  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.660 0.800 2.015 ;
        RECT  0.135 1.660 0.465 2.255 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.909  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 2.480 2.165 3.320 ;
        RECT  1.805 0.535 2.165 3.320 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.940 3.555 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.120 -0.180 1.460 0.505 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.540 0.520 1.430 ;
        RECT  0.180 1.200 1.470 1.430 ;
        RECT  1.160 1.200 1.470 2.860 ;
        RECT  0.180 2.500 1.470 2.860 ;
        RECT  0.180 2.500 0.540 3.335 ;
    END
END CLKBUF_X4_18_SVT_WB

MACRO CLKBUF_X40_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X40_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.548  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.145 0.855 1.685 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.960  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  13.945 0.475 14.305 0.835 ;
        RECT  13.850 1.760 14.235 3.135 ;
        RECT  11.070 0.995 14.235 1.365 ;
        RECT  13.945 0.475 14.235 1.365 ;
        RECT  5.720 1.760 14.235 2.150 ;
        RECT  12.040 0.995 13.060 2.150 ;
        RECT  11.070 0.990 12.860 1.365 ;
        RECT  12.505 0.515 12.860 2.150 ;
        RECT  12.405 0.990 12.775 3.450 ;
        RECT  11.070 0.505 11.425 1.365 ;
        RECT  10.995 1.760 11.345 3.445 ;
        RECT  5.720 0.505 11.425 0.810 ;
        RECT  9.665 1.760 10.025 3.450 ;
        RECT  5.720 0.470 9.955 0.810 ;
        RECT  8.315 1.760 8.715 3.195 ;
        RECT  7.000 1.760 7.405 3.180 ;
        RECT  5.720 0.465 7.315 0.810 ;
        RECT  5.720 1.760 6.040 3.195 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.120 4.100 ;
        RECT  13.150 2.380 13.490 4.100 ;
        RECT  11.710 2.655 12.050 4.100 ;
        RECT  4.990 2.555 5.330 4.100 ;
        RECT  2.220 2.615 2.560 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.120 0.180 ;
        RECT  13.230 -0.180 13.570 0.755 ;
        RECT  11.790 -0.180 12.130 0.760 ;
        RECT  4.990 -0.180 5.330 0.775 ;
        RECT  2.230 -0.180 2.570 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.505 1.865 0.770 ;
        RECT  1.520 0.505 1.865 1.455 ;
        RECT  3.000 0.465 3.235 3.225 ;
        RECT  1.520 1.060 3.235 1.455 ;
        RECT  4.270 0.510 4.610 1.455 ;
        RECT  1.520 1.065 10.435 1.455 ;
        RECT  0.210 2.360 1.820 2.785 ;
        RECT  4.270 0.510 4.565 3.205 ;
        RECT  2.925 1.065 3.260 3.225 ;
        RECT  0.210 2.360 0.540 3.385 ;
        RECT  1.520 0.505 1.820 3.435 ;
        RECT  1.485 2.360 1.820 3.435 ;
    END
END CLKBUF_X40_18_SVT_WB

MACRO CLKBUF_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.340  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.660 0.800 2.015 ;
        RECT  0.135 1.660 0.465 2.255 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.666  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 2.615 2.165 2.935 ;
        RECT  1.805 0.535 2.165 2.935 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.120 -0.180 1.460 0.505 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.540 0.520 1.430 ;
        RECT  0.180 1.200 1.470 1.430 ;
        RECT  1.160 1.200 1.470 2.860 ;
        RECT  0.180 2.500 1.470 2.860 ;
        RECT  0.180 2.500 0.515 3.350 ;
    END
END CLKBUF_X3_18_SVT_WB

MACRO CLKBUF_X32_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X32_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.083  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.705 1.195 2.920 1.755 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.449  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  12.300 1.920 12.640 3.395 ;
        RECT  12.300 0.525 12.640 1.215 ;
        RECT  5.100 1.920 12.640 2.150 ;
        RECT  7.980 0.985 12.640 1.215 ;
        RECT  10.860 1.920 11.200 3.140 ;
        RECT  10.860 0.525 11.200 1.215 ;
        RECT  9.420 1.920 9.760 3.175 ;
        RECT  9.420 0.525 9.760 1.215 ;
        RECT  7.705 0.990 8.610 2.150 ;
        RECT  7.980 0.470 8.320 3.175 ;
        RECT  6.565 0.990 8.610 1.220 ;
        RECT  6.540 1.920 6.880 3.175 ;
        RECT  6.565 0.525 6.880 1.220 ;
        RECT  5.100 0.525 6.880 0.815 ;
        RECT  5.100 1.920 5.440 3.190 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.880 4.100 ;
        RECT  11.580 2.415 11.920 4.100 ;
        RECT  10.140 2.400 10.480 4.100 ;
        RECT  8.700 2.420 9.040 4.100 ;
        RECT  7.260 2.430 7.600 4.100 ;
        RECT  5.820 2.430 6.160 4.100 ;
        RECT  4.340 3.515 4.680 4.100 ;
        RECT  1.500 3.515 1.840 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.880 0.180 ;
        RECT  11.580 -0.180 11.920 0.755 ;
        RECT  10.140 -0.180 10.480 0.755 ;
        RECT  8.700 -0.180 9.040 0.755 ;
        RECT  7.260 -0.180 7.600 0.760 ;
        RECT  4.340 -0.180 4.680 0.405 ;
        RECT  1.500 -0.180 1.840 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.755 0.470 1.075 0.865 ;
        RECT  2.260 0.480 2.610 0.865 ;
        RECT  3.575 0.500 3.920 0.865 ;
        RECT  0.755 0.635 3.920 0.865 ;
        RECT  3.580 0.500 3.920 1.575 ;
        RECT  3.580 1.205 6.335 1.570 ;
        RECT  3.580 1.205 4.870 1.575 ;
        RECT  4.585 1.205 4.870 2.635 ;
        RECT  0.740 2.405 4.870 2.635 ;
        RECT  2.260 2.405 2.600 3.330 ;
        RECT  3.580 2.405 3.920 3.330 ;
        RECT  0.740 2.405 1.080 3.385 ;
    END
END CLKBUF_X32_18_SVT_WB

MACRO CLKBUF_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.304  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.480 0.645 2.390 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.811  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.775 0.470 2.125 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  0.950 3.165 1.290 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  0.950 -0.180 1.290 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.230 0.455 0.470 1.215 ;
        RECT  0.230 0.985 1.440 1.215 ;
        RECT  1.205 0.985 1.440 2.935 ;
        RECT  0.230 2.705 1.440 2.935 ;
        RECT  0.230 2.705 0.570 3.295 ;
    END
END CLKBUF_X2_18_SVT_WB

MACRO CLKBUF_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.514  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.175 0.600 1.760 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.958  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.540 1.990 9.880 3.395 ;
        RECT  4.140 1.990 9.880 2.220 ;
        RECT  7.865 0.985 8.610 2.220 ;
        RECT  8.100 0.525 8.610 2.220 ;
        RECT  8.220 0.525 8.560 3.175 ;
        RECT  5.500 0.985 8.610 1.215 ;
        RECT  6.900 1.990 7.240 3.395 ;
        RECT  6.900 0.525 7.240 1.215 ;
        RECT  5.460 1.990 5.800 3.395 ;
        RECT  5.500 0.525 5.800 1.215 ;
        RECT  4.140 0.525 5.800 0.760 ;
        RECT  4.140 1.990 4.480 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  6.180 2.470 6.520 4.100 ;
        RECT  2.060 3.565 2.400 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  8.940 -0.180 9.280 0.755 ;
        RECT  6.180 -0.180 6.520 0.755 ;
        RECT  0.740 -0.180 1.080 0.770 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.500 0.470 1.840 1.270 ;
        RECT  2.820 0.470 3.160 1.270 ;
        RECT  1.500 1.040 3.910 1.270 ;
        RECT  3.625 1.130 5.190 1.490 ;
        RECT  1.500 2.290 3.910 2.580 ;
        RECT  3.625 1.040 3.910 2.580 ;
        RECT  0.180 2.395 1.840 2.720 ;
        RECT  0.180 2.395 0.520 3.330 ;
        RECT  2.820 2.290 3.160 3.330 ;
    END
END CLKBUF_X24_18_SVT_WB

MACRO CLKBUF_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.283  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.115 0.715 1.660 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.155  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.795 2.430 8.145 3.220 ;
        RECT  5.145 1.085 8.135 1.415 ;
        RECT  7.795 0.525 8.135 1.415 ;
        RECT  6.355 2.430 8.145 2.750 ;
        RECT  6.090 1.085 6.845 2.745 ;
        RECT  6.355 0.525 6.695 3.175 ;
        RECT  5.145 1.080 6.695 1.415 ;
        RECT  3.710 2.430 8.145 2.745 ;
        RECT  5.035 2.430 5.375 3.175 ;
        RECT  5.145 0.525 5.375 1.415 ;
        RECT  3.710 0.525 5.375 0.795 ;
        RECT  3.710 2.430 5.375 2.755 ;
        RECT  3.710 2.430 4.050 3.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.075 3.160 7.415 4.100 ;
        RECT  2.985 3.000 3.330 4.100 ;
        RECT  0.185 2.400 0.525 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.075 -0.180 7.415 0.760 ;
        RECT  2.985 -0.180 3.330 0.790 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.265 0.470 2.605 1.580 ;
        RECT  0.945 0.470 1.285 1.580 ;
        RECT  2.265 1.335 4.815 1.570 ;
        RECT  0.945 1.350 3.480 1.580 ;
        RECT  3.200 1.335 3.480 2.635 ;
        RECT  0.945 2.405 3.480 2.635 ;
        RECT  0.945 2.405 1.285 3.330 ;
        RECT  2.265 2.405 2.605 3.330 ;
    END
END CLKBUF_X20_18_SVT_WB

MACRO CLKBUF_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.969  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.170 1.025 1.730 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.352  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.580 2.150 5.920 3.395 ;
        RECT  2.930 0.985 5.920 1.215 ;
        RECT  5.580 0.525 5.920 1.215 ;
        RECT  4.260 2.150 5.920 2.400 ;
        RECT  4.025 0.985 4.715 2.380 ;
        RECT  4.260 0.525 4.600 3.395 ;
        RECT  2.820 2.150 5.920 2.380 ;
        RECT  2.820 2.150 3.160 3.450 ;
        RECT  2.930 0.465 3.160 1.215 ;
        RECT  2.875 0.465 3.160 0.810 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  3.540 2.610 3.880 4.100 ;
        RECT  0.725 3.565 1.090 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  3.540 -0.180 3.880 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.155 0.510 0.525 0.810 ;
        RECT  1.495 0.515 1.840 0.810 ;
        RECT  0.155 0.580 1.840 0.810 ;
        RECT  1.500 1.445 3.725 1.685 ;
        RECT  0.180 2.575 1.840 2.805 ;
        RECT  0.180 2.575 0.520 2.880 ;
        RECT  1.500 0.515 1.840 3.395 ;
    END
END CLKBUF_X16_18_SVT_WB

MACRO CLKBUF_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKBUF_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.524  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.155 0.710 1.715 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.604  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.075 2.420 5.460 3.470 ;
        RECT  2.260 2.430 5.460 2.740 ;
        RECT  4.040 2.420 5.460 2.740 ;
        RECT  4.040 0.985 4.375 2.740 ;
        RECT  3.700 2.430 4.040 3.175 ;
        RECT  3.700 0.525 4.040 1.215 ;
        RECT  2.260 0.985 4.375 1.215 ;
        RECT  2.260 2.430 2.600 3.395 ;
        RECT  2.260 0.525 2.600 1.215 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  2.980 3.115 3.320 4.100 ;
        RECT  0.180 2.405 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.420 -0.180 4.760 0.755 ;
        RECT  2.980 -0.180 3.320 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 1.485 3.770 1.770 ;
        RECT  0.940 0.590 1.280 3.395 ;
    END
END CLKBUF_X12_18_SVT_WB

MACRO CLKAND2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKAND2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.578  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.425 2.150 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.578  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.605 2.330 2.840 2.560 ;
        RECT  2.500 1.425 2.840 2.560 ;
        RECT  0.605 1.390 0.980 2.560 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.571  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.135 1.200 5.515 2.350 ;
        RECT  3.600 3.130 5.260 3.395 ;
        RECT  4.920 2.120 5.260 3.395 ;
        RECT  3.600 1.200 5.515 1.430 ;
        RECT  3.600 2.675 3.950 3.395 ;
        RECT  3.600 0.920 3.945 1.430 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  5.640 2.695 5.980 4.100 ;
        RECT  1.520 3.515 1.860 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.360 -0.180 4.700 0.875 ;
        RECT  2.720 -0.180 3.060 0.735 ;
        RECT  0.330 -0.180 0.670 0.840 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.595 0.510 1.900 1.195 ;
        RECT  1.595 0.965 3.370 1.195 ;
        RECT  3.070 1.820 4.620 2.160 ;
        RECT  3.070 0.965 3.370 3.170 ;
        RECT  0.760 2.940 3.370 3.170 ;
        RECT  0.760 2.940 1.100 3.385 ;
        RECT  2.280 2.940 2.620 3.450 ;
    END
END CLKAND2_X8_18_SVT_WB

MACRO CLKAND2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKAND2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.125 1.425 1.935 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 2.095 0.530 2.375 ;
        RECT  0.130 1.390 0.470 2.375 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.612  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.860 2.615 4.200 3.330 ;
        RECT  3.165 1.465 3.950 2.955 ;
        RECT  3.165 0.630 3.490 2.955 ;
        RECT  2.420 2.615 4.200 2.955 ;
        RECT  2.420 2.615 2.760 3.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  1.660 3.045 2.000 4.100 ;
        RECT  0.180 2.630 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  2.380 -0.180 2.720 1.385 ;
        RECT  0.190 -0.180 0.530 0.945 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.655 1.780 2.935 2.120 ;
        RECT  1.655 0.605 1.985 2.745 ;
        RECT  0.900 2.405 1.985 2.745 ;
        RECT  0.900 2.405 1.240 3.215 ;
    END
END CLKAND2_X6_18_SVT_WB

MACRO CLKAND2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKAND2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.370 1.315 2.180 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.390 0.470 2.200 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.914  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.150 3.070 1.380 ;
        RECT  2.730 0.870 3.070 1.380 ;
        RECT  2.280 1.150 2.660 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.560 3.125 1.900 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.005 -0.180 2.310 0.920 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.270 0.800 1.775 1.140 ;
        RECT  1.545 1.390 2.050 2.200 ;
        RECT  1.545 0.800 1.775 2.750 ;
        RECT  0.840 2.410 1.775 2.750 ;
        RECT  0.840 2.410 1.180 3.220 ;
    END
END CLKAND2_X4_18_SVT_WB

MACRO CLKAND2_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKAND2_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.390 1.315 2.200 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.288  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.390 0.470 2.200 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.676  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.120 3.070 1.350 ;
        RECT  2.730 0.550 3.070 1.350 ;
        RECT  2.320 1.120 2.660 3.435 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.560 3.110 1.900 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.005 -0.180 2.310 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.270 0.870 1.775 1.160 ;
        RECT  1.545 1.390 2.090 1.780 ;
        RECT  1.545 0.870 1.775 2.770 ;
        RECT  0.840 2.430 1.775 2.770 ;
        RECT  0.840 2.430 1.180 3.230 ;
    END
END CLKAND2_X3_18_SVT_WB

MACRO CLKAND2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKAND2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.820 1.030 2.100 ;
        RECT  0.420 1.535 0.760 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.268  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 1.255 1.590 1.795 ;
        RECT  1.195 1.255 1.590 1.655 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.754  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.795 2.660 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 2.675 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.370 -0.180 1.710 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.795 2.095 1.025 ;
        RECT  0.180 0.795 0.520 1.135 ;
        RECT  1.820 0.795 2.095 2.975 ;
        RECT  0.900 2.635 2.095 2.975 ;
        RECT  0.900 2.635 1.240 3.450 ;
    END
END CLKAND2_X2_18_SVT_WB

MACRO CLKAND2_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKAND2_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.230 1.820 4.320 2.160 ;
        RECT  1.540 2.135 3.570 2.365 ;
        RECT  1.540 1.860 1.880 2.365 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.160 1.360 5.465 1.960 ;
        RECT  0.750 1.360 5.465 1.590 ;
        RECT  2.540 1.360 2.880 1.905 ;
        RECT  0.750 1.360 2.880 1.630 ;
        RECT  0.400 1.805 1.060 2.145 ;
        RECT  0.750 1.360 1.060 2.145 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.206  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.000 0.540 9.340 3.135 ;
        RECT  6.375 1.225 9.340 1.600 ;
        RECT  7.680 0.495 8.020 3.135 ;
        RECT  6.375 1.220 8.020 1.600 ;
        RECT  6.375 0.485 6.700 3.190 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  4.220 3.065 4.560 4.100 ;
        RECT  2.780 3.065 3.120 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  5.450 -0.180 5.890 0.410 ;
        RECT  2.740 -0.180 3.080 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.340 0.640 6.025 0.980 ;
        RECT  5.795 1.020 6.145 1.425 ;
        RECT  5.795 0.640 6.025 2.825 ;
        RECT  0.740 2.595 6.025 2.825 ;
        RECT  2.060 2.595 3.840 2.835 ;
        RECT  2.060 2.595 2.400 3.405 ;
        RECT  3.500 2.595 3.840 3.405 ;
        RECT  4.925 2.595 5.280 3.405 ;
        RECT  0.740 2.595 1.075 3.445 ;
    END
END CLKAND2_X16_18_SVT_WB

MACRO CLKAND2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN CLKAND2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.578  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.430 1.445 2.240 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.578  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.640 2.330 2.960 2.670 ;
        RECT  2.620 1.445 2.960 2.670 ;
        RECT  0.640 1.390 0.980 2.670 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.614  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.675 2.170 7.015 3.335 ;
        RECT  3.790 2.170 7.015 2.425 ;
        RECT  5.180 2.170 5.575 3.395 ;
        RECT  5.235 0.585 5.575 3.395 ;
        RECT  3.795 0.590 5.575 0.930 ;
        RECT  5.180 0.585 5.575 0.930 ;
        RECT  3.795 2.170 4.135 3.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  5.955 2.655 6.295 4.100 ;
        RECT  4.515 2.655 4.855 4.100 ;
        RECT  1.620 3.515 1.960 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  5.995 -0.180 6.340 0.890 ;
        RECT  3.035 -0.180 3.375 0.755 ;
        RECT  0.430 -0.180 0.770 0.945 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.660 0.605 2.000 1.215 ;
        RECT  1.660 0.985 3.560 1.215 ;
        RECT  3.330 1.170 4.365 1.510 ;
        RECT  3.330 0.985 3.560 3.170 ;
        RECT  0.860 2.940 3.560 3.170 ;
        RECT  0.860 2.940 1.200 3.385 ;
        RECT  2.380 2.940 2.720 3.450 ;
    END
END CLKAND2_X12_18_SVT_WB

MACRO BUF_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.671  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 1.750 0.860 2.175 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.385 2.545 3.725 3.385 ;
        RECT  2.065 1.055 3.725 1.350 ;
        RECT  3.385 0.535 3.725 1.350 ;
        RECT  2.065 2.545 3.725 2.940 ;
        RECT  2.860 1.055 3.235 2.940 ;
        RECT  2.065 0.590 2.415 1.350 ;
        RECT  2.065 2.545 2.405 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  1.300 3.570 1.640 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  1.300 -0.180 1.640 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.905 1.425 1.160 ;
        RECT  1.090 0.905 1.425 2.670 ;
        RECT  1.090 1.620 2.605 1.960 ;
        RECT  1.090 1.620 1.430 2.670 ;
        RECT  0.740 2.405 1.430 2.670 ;
    END
END BUF_X8_18_SVT_WB

MACRO BUF_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.274  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.665 0.600 2.175 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.820 2.585 3.160 3.390 ;
        RECT  1.500 1.110 3.160 1.435 ;
        RECT  2.820 0.615 3.160 1.435 ;
        RECT  1.500 2.585 3.160 2.920 ;
        RECT  2.370 1.110 2.715 2.920 ;
        RECT  1.500 0.615 1.870 1.435 ;
        RECT  1.500 2.585 1.850 3.395 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.730 3.555 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.740 -0.180 1.080 0.360 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 1.125 1.365 ;
        RECT  0.830 1.665 2.140 1.960 ;
        RECT  0.830 1.100 1.125 2.690 ;
        RECT  0.170 2.450 1.125 2.690 ;
    END
END BUF_X6_18_SVT_WB

MACRO BUF_X5_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X5_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.750 0.755 2.180 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.718  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.500 2.380 3.160 2.790 ;
        RECT  1.500 1.010 3.160 1.340 ;
        RECT  2.345 1.010 2.720 2.790 ;
        RECT  1.500 2.380 1.855 3.310 ;
        RECT  1.500 0.535 1.840 1.340 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.255 3.425 2.605 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.260 -0.180 2.600 0.490 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.535 0.520 1.440 ;
        RECT  0.180 1.105 1.270 1.440 ;
        RECT  1.040 1.620 1.610 1.960 ;
        RECT  1.040 1.105 1.270 2.750 ;
        RECT  0.180 2.410 1.270 2.750 ;
        RECT  0.180 2.410 0.520 3.220 ;
    END
END BUF_X5_18_SVT_WB

MACRO BUF_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.720 1.010 2.180 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.535 2.135 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.940 -0.180 1.280 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.535 0.520 1.485 ;
        RECT  0.180 1.255 1.470 1.485 ;
        RECT  1.240 1.255 1.470 2.750 ;
        RECT  0.180 2.410 1.470 2.750 ;
        RECT  0.180 2.410 0.520 3.385 ;
    END
END BUF_X4_18_SVT_WB

MACRO BUF_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.296  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.660 0.800 2.015 ;
        RECT  0.135 1.660 0.465 2.255 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.888  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.700 0.760 2.110 2.935 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  0.940 -0.180 1.280 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.905 0.520 1.430 ;
        RECT  0.180 1.200 1.470 1.430 ;
        RECT  1.160 1.200 1.470 3.130 ;
        RECT  0.180 2.770 1.470 3.130 ;
    END
END BUF_X3_18_SVT_WB

MACRO BUF_X32_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X32_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 2.111  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.130 1.705 3.150 2.265 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 9.504  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.420 2.550 14.760 3.285 ;
        RECT  4.790 1.110 14.760 1.360 ;
        RECT  14.420 0.585 14.760 1.360 ;
        RECT  4.840 2.550 14.760 2.890 ;
        RECT  13.100 2.550 13.440 3.290 ;
        RECT  13.100 0.585 13.440 1.360 ;
        RECT  11.775 2.550 12.120 3.290 ;
        RECT  11.775 0.585 12.120 1.360 ;
        RECT  10.340 2.550 10.680 3.390 ;
        RECT  10.340 0.585 10.680 1.360 ;
        RECT  10.080 1.110 10.540 2.890 ;
        RECT  9.020 2.550 9.360 3.390 ;
        RECT  9.020 0.585 9.360 1.360 ;
        RECT  7.580 2.550 7.920 3.390 ;
        RECT  7.580 0.585 7.920 1.360 ;
        RECT  6.260 2.550 6.600 3.390 ;
        RECT  6.260 0.585 6.600 1.360 ;
        RECT  4.840 2.550 5.160 3.390 ;
        RECT  4.790 0.585 5.160 1.360 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.680 4.100 ;
        RECT  15.140 2.640 15.480 4.100 ;
        RECT  11.060 3.160 11.400 4.100 ;
        RECT  8.300 3.160 8.640 4.100 ;
        RECT  5.540 3.155 5.880 4.100 ;
        RECT  1.460 3.150 1.800 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.680 0.180 ;
        RECT  15.140 -0.180 15.480 1.395 ;
        RECT  11.060 -0.180 11.400 0.760 ;
        RECT  8.300 -0.180 8.640 0.760 ;
        RECT  5.540 -0.180 5.880 0.765 ;
        RECT  1.460 -0.180 1.800 0.925 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.585 1.080 1.395 ;
        RECT  2.180 0.585 2.520 1.395 ;
        RECT  0.740 1.165 3.840 1.395 ;
        RECT  3.500 1.625 9.655 1.965 ;
        RECT  0.740 2.610 3.840 2.885 ;
        RECT  3.500 0.585 3.840 3.390 ;
        RECT  0.740 2.610 1.075 3.405 ;
        RECT  2.180 2.610 2.520 3.450 ;
    END
END BUF_X32_18_SVT_WB

MACRO BUF_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.525 1.705 0.980 2.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 0.470 2.100 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.240 4.100 ;
        RECT  1.000 3.165 1.340 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.240 0.180 ;
        RECT  1.000 -0.180 1.340 0.755 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.280 0.575 0.620 1.215 ;
        RECT  0.280 0.985 1.490 1.215 ;
        RECT  1.210 0.985 1.490 2.935 ;
        RECT  0.280 2.705 1.490 2.935 ;
        RECT  0.280 2.705 0.620 3.295 ;
    END
END BUF_X2_18_SVT_WB

MACRO BUF_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.635 1.915 2.230 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 7.128  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  11.020 2.525 11.360 3.385 ;
        RECT  3.940 1.030 11.360 1.320 ;
        RECT  11.020 0.470 11.360 1.320 ;
        RECT  3.940 2.525 11.360 2.865 ;
        RECT  9.700 2.525 10.040 3.385 ;
        RECT  9.700 0.470 10.040 1.320 ;
        RECT  8.260 2.525 8.600 3.385 ;
        RECT  8.260 0.470 8.600 1.320 ;
        RECT  7.955 1.030 8.380 2.865 ;
        RECT  6.820 2.525 7.160 3.385 ;
        RECT  6.820 0.470 7.160 1.320 ;
        RECT  5.380 2.525 5.720 3.385 ;
        RECT  5.380 0.470 5.720 1.320 ;
        RECT  3.940 2.525 4.280 3.385 ;
        RECT  3.940 0.535 4.280 1.320 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 12.320 4.100 ;
        RECT  11.740 2.575 12.080 4.100 ;
        RECT  8.980 3.135 9.320 4.100 ;
        RECT  7.540 3.145 7.880 4.100 ;
        RECT  6.100 3.095 6.440 4.100 ;
        RECT  4.660 3.095 5.000 4.100 ;
        RECT  3.180 3.005 3.520 4.100 ;
        RECT  1.660 3.515 2.000 4.100 ;
        RECT  0.180 2.625 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 12.320 0.180 ;
        RECT  11.740 -0.180 12.080 1.280 ;
        RECT  8.980 -0.180 9.320 0.760 ;
        RECT  7.540 -0.180 7.880 0.760 ;
        RECT  6.100 -0.180 6.440 0.760 ;
        RECT  4.660 -0.180 5.000 0.760 ;
        RECT  3.180 -0.180 3.520 0.875 ;
        RECT  1.660 -0.180 2.000 0.875 ;
        RECT  0.180 -0.180 0.520 1.345 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 0.535 1.240 1.345 ;
        RECT  0.900 1.115 2.760 1.345 ;
        RECT  2.420 1.620 7.360 1.960 ;
        RECT  0.900 2.520 2.760 2.810 ;
        RECT  0.900 2.520 1.240 3.280 ;
        RECT  2.420 0.535 2.760 3.385 ;
    END
END BUF_X24_18_SVT_WB

MACRO BUF_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.550 1.665 1.135 2.210 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.940  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.940 2.465 9.280 3.390 ;
        RECT  3.540 0.990 9.280 1.265 ;
        RECT  8.940 0.470 9.280 1.265 ;
        RECT  7.620 2.465 9.280 2.810 ;
        RECT  7.620 2.465 7.960 3.390 ;
        RECT  7.620 0.470 7.960 1.265 ;
        RECT  6.300 2.465 9.280 2.805 ;
        RECT  6.300 0.470 6.640 3.390 ;
        RECT  3.540 2.475 6.640 2.815 ;
        RECT  4.860 2.475 5.200 3.390 ;
        RECT  3.540 0.985 5.200 1.265 ;
        RECT  4.860 0.470 5.200 1.265 ;
        RECT  3.540 2.475 3.880 3.390 ;
        RECT  3.540 0.470 3.880 1.265 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  5.580 3.160 5.920 4.100 ;
        RECT  0.180 2.580 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  5.580 -0.180 5.920 0.760 ;
        RECT  0.180 -0.180 0.520 1.275 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.885 0.540 1.260 1.375 ;
        RECT  0.885 1.135 2.560 1.375 ;
        RECT  2.220 1.620 5.870 1.960 ;
        RECT  0.900 2.620 2.560 2.850 ;
        RECT  0.900 2.620 1.240 3.390 ;
        RECT  2.220 0.540 2.560 3.390 ;
    END
END BUF_X20_18_SVT_WB

MACRO BUF_X18_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X18_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.675 1.690 1.485 2.225 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.808  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.995 2.555 9.335 3.385 ;
        RECT  3.235 0.995 9.335 1.350 ;
        RECT  8.995 0.470 9.335 1.350 ;
        RECT  3.235 2.560 9.335 2.875 ;
        RECT  6.265 2.555 9.335 2.875 ;
        RECT  7.555 2.555 7.895 3.385 ;
        RECT  7.555 0.470 7.895 1.350 ;
        RECT  6.265 0.995 6.910 2.875 ;
        RECT  6.115 2.560 6.455 3.385 ;
        RECT  6.115 0.535 6.455 1.350 ;
        RECT  4.675 2.560 5.015 3.385 ;
        RECT  4.675 0.535 5.015 1.350 ;
        RECT  3.235 2.560 3.575 3.385 ;
        RECT  3.235 0.535 3.575 1.350 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  8.275 3.155 8.615 4.100 ;
        RECT  6.835 3.160 7.175 4.100 ;
        RECT  5.395 3.155 5.735 4.100 ;
        RECT  3.955 3.160 4.295 4.100 ;
        RECT  2.475 3.050 2.815 4.100 ;
        RECT  0.955 3.515 1.295 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  8.275 -0.180 8.615 0.765 ;
        RECT  6.835 -0.180 7.175 0.765 ;
        RECT  5.395 -0.180 5.735 0.765 ;
        RECT  3.955 -0.180 4.295 0.765 ;
        RECT  2.475 -0.180 2.815 0.875 ;
        RECT  0.955 -0.180 1.295 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.195 0.535 0.535 1.345 ;
        RECT  0.195 1.105 2.055 1.345 ;
        RECT  1.715 1.620 6.035 1.960 ;
        RECT  0.195 2.570 2.055 2.875 ;
        RECT  0.195 2.570 0.535 3.385 ;
        RECT  1.715 0.535 2.055 3.385 ;
    END
END BUF_X18_18_SVT_WB

MACRO BUF_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.515 1.760 1.780 2.100 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.752  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.660 2.420 8.000 3.230 ;
        RECT  3.580 1.050 8.000 1.390 ;
        RECT  7.660 0.580 8.000 1.390 ;
        RECT  3.580 2.420 8.000 2.760 ;
        RECT  6.340 2.420 6.680 3.230 ;
        RECT  6.340 0.580 6.680 1.390 ;
        RECT  6.235 1.050 6.595 2.760 ;
        RECT  5.020 2.420 5.360 3.230 ;
        RECT  5.020 0.580 5.360 1.390 ;
        RECT  3.580 2.420 3.920 3.230 ;
        RECT  3.580 0.590 3.920 1.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  8.380 2.420 8.720 4.100 ;
        RECT  4.300 3.110 4.640 4.100 ;
        RECT  1.500 3.515 1.840 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.380 -0.180 8.720 1.390 ;
        RECT  4.300 -0.180 4.640 0.810 ;
        RECT  1.500 -0.180 1.840 0.970 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.740 0.535 1.080 1.440 ;
        RECT  0.740 1.200 2.600 1.440 ;
        RECT  2.260 1.620 6.005 1.960 ;
        RECT  0.740 2.380 2.600 2.720 ;
        RECT  0.740 2.380 1.080 3.385 ;
        RECT  2.260 0.535 2.600 3.385 ;
    END
END BUF_X16_18_SVT_WB

MACRO BUF_X14_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X14_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.923  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.255 1.480 1.725 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.620  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.280 2.375 7.620 3.390 ;
        RECT  3.080 0.995 7.620 1.295 ;
        RECT  7.280 0.465 7.620 1.295 ;
        RECT  3.080 2.375 7.620 2.730 ;
        RECT  5.840 2.375 6.180 3.245 ;
        RECT  5.840 0.470 6.180 1.295 ;
        RECT  5.140 0.995 5.505 2.730 ;
        RECT  4.520 2.375 4.860 3.225 ;
        RECT  4.520 0.470 4.860 1.295 ;
        RECT  3.080 2.375 4.860 2.735 ;
        RECT  3.080 2.375 3.420 3.225 ;
        RECT  3.080 0.470 3.420 1.295 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  6.560 3.100 6.900 4.100 ;
        RECT  3.800 3.145 4.140 4.100 ;
        RECT  1.040 2.635 1.380 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  6.560 -0.180 6.900 0.765 ;
        RECT  3.800 -0.180 4.140 0.765 ;
        RECT  1.000 -0.180 1.340 0.410 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.240 0.540 0.580 0.920 ;
        RECT  0.240 0.690 2.100 0.920 ;
        RECT  1.760 1.620 4.690 1.960 ;
        RECT  0.265 2.065 2.100 2.405 ;
        RECT  0.265 2.065 0.545 3.445 ;
        RECT  1.760 0.690 2.100 3.445 ;
    END
END BUF_X14_18_SVT_WB

MACRO BUF_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.660 0.710 2.225 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.020 2.450 5.360 3.385 ;
        RECT  2.260 1.105 5.360 1.345 ;
        RECT  5.020 0.535 5.360 1.345 ;
        RECT  2.260 2.450 5.360 2.755 ;
        RECT  4.020 1.105 4.405 2.755 ;
        RECT  3.700 2.450 4.040 3.385 ;
        RECT  3.700 0.535 4.040 1.345 ;
        RECT  2.260 2.450 2.600 3.385 ;
        RECT  2.260 0.535 2.600 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  2.980 3.070 3.320 4.100 ;
        RECT  0.165 2.545 0.535 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  2.980 -0.180 3.320 0.855 ;
        RECT  0.180 -0.180 0.520 1.345 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.940 0.535 1.275 3.385 ;
        RECT  0.940 1.620 3.790 1.960 ;
        RECT  0.940 1.425 1.280 3.385 ;
    END
END BUF_X12_18_SVT_WB

MACRO BUF_X10_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUF_X10_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.595 1.770 1.200 2.150 ;
        END
    END A
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.432  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.065 2.610 5.405 3.390 ;
        RECT  2.305 0.990 5.405 1.275 ;
        RECT  5.065 0.470 5.405 1.275 ;
        RECT  2.305 2.610 5.405 2.885 ;
        RECT  3.625 2.610 3.965 3.390 ;
        RECT  3.625 0.470 3.965 1.275 ;
        RECT  3.380 0.990 3.790 2.885 ;
        RECT  2.305 2.610 2.645 3.430 ;
        RECT  2.305 0.470 2.645 1.275 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.345 3.160 4.685 4.100 ;
        RECT  0.240 2.575 0.580 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.345 -0.180 4.685 0.760 ;
        RECT  0.240 -0.180 0.580 1.360 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.975 0.475 1.315 1.295 ;
        RECT  0.975 1.010 1.910 1.295 ;
        RECT  1.550 1.010 1.910 1.960 ;
        RECT  1.550 1.620 2.880 1.960 ;
        RECT  1.550 1.010 1.905 2.930 ;
        RECT  0.975 2.565 1.905 2.930 ;
        RECT  0.975 2.565 1.300 3.385 ;
    END
END BUF_X10_18_SVT_WB

MACRO BUFT_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.264  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.125 1.905 3.580 2.295 ;
        RECT  2.690 1.820 3.375 2.140 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.540 0.835 1.885 ;
        RECT  0.140 1.540 0.455 2.160 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.197  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.775 3.080 6.580 3.425 ;
        RECT  6.255 0.520 6.580 3.425 ;
        RECT  5.990 2.585 6.580 3.425 ;
        RECT  4.525 0.520 6.580 0.755 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  6.810 2.610 7.050 4.100 ;
        RECT  3.235 3.570 3.600 4.100 ;
        RECT  0.860 3.430 1.225 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.810 -0.180 7.055 1.265 ;
        RECT  3.765 -0.180 4.105 0.350 ;
        RECT  0.765 -0.180 0.995 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.260 0.410 1.605 0.895 ;
        RECT  0.180 0.895 1.310 1.125 ;
        RECT  0.180 0.845 0.465 1.175 ;
        RECT  1.080 0.665 1.310 2.620 ;
        RECT  1.080 2.165 2.460 2.400 ;
        RECT  0.235 2.390 1.330 2.620 ;
        RECT  0.235 2.390 0.465 2.825 ;
        RECT  2.325 1.155 2.625 1.590 ;
        RECT  2.325 1.360 3.835 1.590 ;
        RECT  3.605 1.445 4.085 1.675 ;
        RECT  3.810 1.955 4.500 2.305 ;
        RECT  2.690 2.525 4.085 2.765 ;
        RECT  3.810 1.445 4.085 2.765 ;
        RECT  1.640 2.630 2.920 2.860 ;
        RECT  1.640 2.630 1.980 3.035 ;
        RECT  1.835 0.655 3.400 0.885 ;
        RECT  3.060 0.855 4.295 1.095 ;
        RECT  4.065 0.985 5.665 1.215 ;
        RECT  1.835 0.655 2.065 1.450 ;
        RECT  1.540 1.190 2.065 1.450 ;
        RECT  5.395 0.985 5.665 1.860 ;
        RECT  4.800 1.540 5.665 1.860 ;
        RECT  4.800 1.540 5.045 2.765 ;
        RECT  4.315 2.535 5.045 2.765 ;
        RECT  4.315 2.535 4.545 3.320 ;
        RECT  2.360 3.090 4.545 3.320 ;
    END
END BUFT_X8_18_SVT_WB

MACRO BUFT_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.264  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.395 1.905 3.740 2.295 ;
        RECT  2.850 1.905 3.740 2.160 ;
        RECT  2.850 1.820 3.335 2.160 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.466  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.545 1.540 0.995 2.160 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.077  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.275 0.520 6.580 3.080 ;
        RECT  4.935 3.080 6.560 3.420 ;
        RECT  4.675 0.520 6.580 0.755 ;
        RECT  4.935 3.080 5.165 3.470 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  3.395 3.570 3.760 4.100 ;
        RECT  1.020 3.430 1.385 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  3.925 -0.180 4.265 0.350 ;
        RECT  0.925 -0.180 1.155 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.420 0.410 1.765 0.895 ;
        RECT  0.340 0.895 1.470 1.125 ;
        RECT  0.340 0.845 0.625 1.175 ;
        RECT  1.240 0.665 1.470 2.620 ;
        RECT  1.240 2.165 2.620 2.400 ;
        RECT  0.395 2.390 1.490 2.620 ;
        RECT  0.395 2.390 0.625 2.825 ;
        RECT  2.485 1.155 2.785 1.590 ;
        RECT  2.485 1.360 3.820 1.590 ;
        RECT  3.565 1.445 4.245 1.675 ;
        RECT  3.970 1.955 4.660 2.305 ;
        RECT  2.850 2.525 4.245 2.765 ;
        RECT  3.970 1.445 4.245 2.765 ;
        RECT  1.800 2.630 3.080 2.860 ;
        RECT  1.800 2.630 2.140 3.035 ;
        RECT  1.995 0.655 3.595 0.885 ;
        RECT  3.175 0.750 4.325 1.095 ;
        RECT  4.050 0.985 5.825 1.215 ;
        RECT  1.995 0.655 2.225 1.450 ;
        RECT  1.700 1.190 2.225 1.450 ;
        RECT  5.555 0.985 5.825 1.860 ;
        RECT  4.960 1.540 5.825 1.860 ;
        RECT  4.960 1.540 5.205 2.765 ;
        RECT  4.475 2.535 5.205 2.765 ;
        RECT  4.475 2.535 4.705 3.320 ;
        RECT  2.520 3.090 4.705 3.320 ;
    END
END BUFT_X6_18_SVT_WB

MACRO BUFT_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.070 3.260 1.720 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.320  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.145 1.015 1.840 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.080  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.960 2.640 4.340 3.430 ;
        RECT  4.110 1.055 4.340 3.430 ;
        RECT  3.960 1.055 4.340 1.710 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  1.035 -0.180 1.375 0.805 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.510 0.655 0.800 ;
        RECT  0.115 0.510 0.345 3.450 ;
        RECT  1.275 1.080 1.615 2.470 ;
        RECT  0.115 2.130 1.615 2.470 ;
        RECT  0.115 2.130 0.430 3.450 ;
        RECT  0.115 3.115 0.520 3.450 ;
        RECT  2.405 1.170 2.640 2.180 ;
        RECT  2.405 1.950 2.965 2.180 ;
        RECT  3.420 1.960 3.855 2.385 ;
        RECT  2.735 1.950 2.965 3.450 ;
        RECT  2.545 3.110 2.965 3.450 ;
        RECT  3.420 1.960 3.715 3.450 ;
        RECT  2.545 3.175 3.715 3.450 ;
        RECT  1.945 0.520 3.355 0.825 ;
        RECT  1.945 0.595 4.805 0.825 ;
        RECT  4.570 0.595 4.805 1.870 ;
        RECT  1.945 0.520 2.175 2.805 ;
        RECT  1.945 2.410 2.505 2.805 ;
    END
END BUFT_X4_18_SVT_WB

MACRO BUFT_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.070 3.260 1.720 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.145 1.015 1.840 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.710  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.960 2.640 4.340 2.930 ;
        RECT  4.110 1.055 4.340 2.930 ;
        RECT  3.960 1.055 4.340 1.710 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.520 3.550 4.865 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.510 -0.180 4.870 0.350 ;
        RECT  1.035 -0.180 1.375 0.805 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.510 0.655 0.800 ;
        RECT  0.115 0.510 0.345 3.450 ;
        RECT  1.275 1.080 1.615 2.470 ;
        RECT  0.115 2.130 1.615 2.470 ;
        RECT  0.115 2.130 0.430 3.450 ;
        RECT  0.115 3.115 0.520 3.450 ;
        RECT  2.405 1.170 2.640 2.180 ;
        RECT  2.405 1.950 2.965 2.180 ;
        RECT  3.420 1.960 3.855 2.385 ;
        RECT  2.735 1.950 2.965 3.450 ;
        RECT  2.545 3.110 2.965 3.450 ;
        RECT  3.420 1.960 3.715 3.450 ;
        RECT  2.545 3.175 3.715 3.450 ;
        RECT  1.945 0.520 3.355 0.825 ;
        RECT  1.945 0.595 4.805 0.825 ;
        RECT  4.570 0.595 4.805 1.870 ;
        RECT  1.945 0.520 2.175 2.805 ;
        RECT  1.945 2.410 2.505 2.805 ;
    END
END BUFT_X3_18_SVT_WB

MACRO BUFT_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.870 1.070 3.260 1.720 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.145 1.015 1.840 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.631  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.960 0.960 4.340 2.930 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  1.035 -0.180 1.375 0.805 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.115 0.510 0.655 0.800 ;
        RECT  0.115 0.510 0.345 3.450 ;
        RECT  1.275 1.080 1.615 2.470 ;
        RECT  0.115 2.130 1.615 2.470 ;
        RECT  0.115 2.130 0.430 3.450 ;
        RECT  0.115 3.115 0.520 3.450 ;
        RECT  2.405 1.170 2.640 2.180 ;
        RECT  2.405 1.950 2.965 2.180 ;
        RECT  2.735 1.950 2.965 3.450 ;
        RECT  2.545 3.110 2.965 3.450 ;
        RECT  2.545 3.175 4.070 3.450 ;
        RECT  3.740 3.175 4.070 3.510 ;
        RECT  3.495 0.410 4.080 0.695 ;
        RECT  1.945 0.520 3.665 0.770 ;
        RECT  1.945 0.520 2.175 2.805 ;
        RECT  1.945 2.410 2.505 2.805 ;
    END
END BUFT_X2_18_SVT_WB

MACRO BUFT_X24_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X24_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.362  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.200 1.975 6.540 2.420 ;
        RECT  5.555 1.785 6.190 2.420 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.126  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.950 0.850 2.365 ;
        RECT  0.140 1.690 0.435 2.365 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 6.042  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  15.380 2.580 15.710 3.340 ;
        RECT  8.665 1.050 15.635 1.280 ;
        RECT  15.380 0.450 15.635 1.280 ;
        RECT  8.625 2.580 15.710 2.815 ;
        RECT  14.050 2.580 14.380 3.340 ;
        RECT  14.070 0.470 14.310 1.280 ;
        RECT  8.625 2.580 14.380 2.820 ;
        RECT  13.565 1.050 13.930 2.820 ;
        RECT  8.665 1.050 13.930 1.290 ;
        RECT  12.650 2.580 12.890 3.340 ;
        RECT  12.630 0.470 12.870 1.290 ;
        RECT  8.625 2.580 12.890 2.825 ;
        RECT  11.325 2.580 11.570 3.340 ;
        RECT  11.305 0.470 11.550 1.290 ;
        RECT  10.010 2.580 10.250 3.365 ;
        RECT  9.990 0.470 10.230 1.290 ;
        RECT  8.625 2.580 8.930 3.340 ;
        RECT  8.665 0.480 8.910 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 16.240 4.100 ;
        RECT  13.375 3.105 13.605 4.100 ;
        RECT  7.820 3.570 8.220 4.100 ;
        RECT  0.890 3.515 1.125 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 16.240 0.180 ;
        RECT  13.300 -0.180 13.640 0.755 ;
        RECT  7.915 -0.180 8.145 0.405 ;
        RECT  0.795 -0.180 1.025 0.425 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.270 0.410 1.610 0.640 ;
        RECT  0.160 0.945 1.500 1.200 ;
        RECT  1.270 0.410 1.500 1.575 ;
        RECT  1.190 2.130 2.740 2.370 ;
        RECT  1.190 0.945 1.420 2.935 ;
        RECT  0.175 2.640 1.420 2.935 ;
        RECT  3.915 1.160 7.060 1.390 ;
        RECT  6.830 1.160 7.060 1.770 ;
        RECT  2.480 1.160 2.835 1.795 ;
        RECT  6.830 1.495 7.860 1.770 ;
        RECT  3.915 1.160 4.205 1.795 ;
        RECT  2.480 1.565 4.205 1.795 ;
        RECT  7.545 1.495 7.860 2.880 ;
        RECT  1.650 2.650 7.860 2.880 ;
        RECT  1.650 2.650 1.965 3.005 ;
        RECT  2.000 0.700 8.395 0.930 ;
        RECT  7.290 0.700 7.685 1.150 ;
        RECT  1.735 0.920 2.250 1.225 ;
        RECT  3.180 0.700 3.560 1.225 ;
        RECT  8.165 1.525 13.155 1.765 ;
        RECT  8.165 0.700 8.395 3.340 ;
        RECT  2.375 3.110 8.395 3.340 ;
        RECT  2.375 3.110 2.665 3.390 ;
        RECT  3.955 3.110 4.185 3.390 ;
    END
END BUFT_X24_18_SVT_WB

MACRO BUFT_X20_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X20_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.986  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.200 1.975 6.540 2.420 ;
        RECT  5.555 1.785 6.190 2.420 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.796  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.950 0.850 2.365 ;
        RECT  0.140 1.690 0.435 2.365 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 5.130  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  14.050 2.580 14.395 3.340 ;
        RECT  8.665 1.050 14.310 1.280 ;
        RECT  14.070 0.470 14.310 1.280 ;
        RECT  8.625 2.580 14.395 2.820 ;
        RECT  12.650 2.580 12.890 3.340 ;
        RECT  12.630 0.470 12.870 1.280 ;
        RECT  12.405 1.050 12.770 2.825 ;
        RECT  8.625 2.580 12.890 2.825 ;
        RECT  8.665 1.050 12.770 1.290 ;
        RECT  11.325 2.580 11.570 3.340 ;
        RECT  11.305 0.470 11.550 1.290 ;
        RECT  10.010 2.580 10.250 3.365 ;
        RECT  9.990 0.470 10.230 1.290 ;
        RECT  8.625 2.580 8.930 3.340 ;
        RECT  8.665 0.480 8.910 1.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 15.120 4.100 ;
        RECT  13.375 3.105 13.605 4.100 ;
        RECT  7.820 3.570 8.220 4.100 ;
        RECT  0.890 3.515 1.125 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 15.120 0.180 ;
        RECT  13.300 -0.180 13.640 0.755 ;
        RECT  7.915 -0.180 8.145 0.405 ;
        RECT  0.795 -0.180 1.025 0.425 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.270 0.410 1.610 0.640 ;
        RECT  0.160 0.945 1.500 1.200 ;
        RECT  1.270 0.410 1.500 1.575 ;
        RECT  1.190 2.130 2.740 2.370 ;
        RECT  1.190 0.945 1.420 2.935 ;
        RECT  0.175 2.640 1.420 2.935 ;
        RECT  3.915 1.160 7.060 1.390 ;
        RECT  6.830 1.160 7.060 1.770 ;
        RECT  2.480 1.160 2.835 1.795 ;
        RECT  6.830 1.495 7.860 1.770 ;
        RECT  3.915 1.160 4.205 1.795 ;
        RECT  2.480 1.565 4.205 1.795 ;
        RECT  7.545 1.495 7.860 2.880 ;
        RECT  1.650 2.650 7.860 2.880 ;
        RECT  1.650 2.650 1.965 3.005 ;
        RECT  2.000 0.700 8.395 0.930 ;
        RECT  7.290 0.700 7.680 1.150 ;
        RECT  1.735 0.920 2.250 1.225 ;
        RECT  3.180 0.700 3.560 1.225 ;
        RECT  8.165 1.525 11.760 1.765 ;
        RECT  8.165 0.700 8.395 3.340 ;
        RECT  2.375 3.110 8.395 3.340 ;
        RECT  2.375 3.110 2.665 3.390 ;
        RECT  3.955 3.110 4.185 3.390 ;
    END
END BUFT_X20_18_SVT_WB

MACRO BUFT_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.400 1.705 3.830 2.205 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.302  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.145 1.015 1.840 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.960 3.010 4.340 3.295 ;
        RECT  4.065 0.510 4.340 3.295 ;
        RECT  4.060 1.705 4.340 2.200 ;
        RECT  3.935 0.510 4.340 0.840 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  1.035 -0.180 1.375 0.805 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.140 0.510 0.655 0.800 ;
        RECT  0.140 0.510 0.370 3.450 ;
        RECT  1.275 1.080 1.615 2.470 ;
        RECT  0.140 2.130 1.615 2.470 ;
        RECT  0.140 2.130 0.430 3.450 ;
        RECT  0.140 3.115 0.520 3.450 ;
        RECT  2.515 1.170 2.805 2.180 ;
        RECT  2.515 1.910 3.170 2.180 ;
        RECT  2.940 1.910 3.170 3.450 ;
        RECT  3.575 2.435 3.835 2.775 ;
        RECT  2.940 2.490 3.835 2.775 ;
        RECT  2.940 2.490 3.245 3.450 ;
        RECT  2.545 3.110 3.245 3.450 ;
        RECT  1.945 0.520 3.600 0.860 ;
        RECT  3.370 0.520 3.600 1.475 ;
        RECT  3.370 1.095 3.835 1.475 ;
        RECT  1.945 0.520 2.285 1.560 ;
        RECT  1.845 1.170 2.285 1.560 ;
        RECT  2.055 0.520 2.285 2.760 ;
        RECT  2.055 2.410 2.595 2.760 ;
    END
END BUFT_X1_18_SVT_WB

MACRO BUFT_X16_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X16_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.878  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.210 1.735 3.890 2.270 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.656  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.735 0.790 2.415 ;
        RECT  0.140 1.735 0.790 2.150 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.320  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.505 2.530 10.290 2.770 ;
        RECT  9.980 0.470 10.290 1.285 ;
        RECT  8.505 2.525 9.995 2.770 ;
        RECT  9.340 1.000 9.995 2.770 ;
        RECT  5.830 1.000 10.290 1.230 ;
        RECT  5.910 3.160 8.840 3.450 ;
        RECT  8.505 2.525 8.840 3.450 ;
        RECT  8.480 0.470 8.825 1.230 ;
        RECT  5.910 3.080 7.535 3.450 ;
        RECT  7.165 0.530 7.515 1.230 ;
        RECT  5.830 0.480 6.185 1.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  10.655 2.665 11.000 4.100 ;
        RECT  9.215 3.060 9.555 4.100 ;
        RECT  3.765 3.570 4.105 4.100 ;
        RECT  0.795 3.515 1.025 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  10.645 -0.180 11.000 1.270 ;
        RECT  9.205 -0.180 9.545 0.755 ;
        RECT  3.765 -0.180 4.105 0.350 ;
        RECT  0.795 -0.180 1.025 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.260 0.410 1.600 0.640 ;
        RECT  1.030 0.635 1.490 0.865 ;
        RECT  0.180 0.985 1.260 1.235 ;
        RECT  0.180 0.920 0.465 1.300 ;
        RECT  1.030 0.635 1.260 1.840 ;
        RECT  1.095 1.615 1.385 2.475 ;
        RECT  1.095 2.195 2.620 2.475 ;
        RECT  0.190 2.730 0.475 3.120 ;
        RECT  1.095 1.615 1.325 3.120 ;
        RECT  0.190 2.890 1.325 3.120 ;
        RECT  2.400 1.165 4.350 1.505 ;
        RECT  4.120 1.165 4.350 2.285 ;
        RECT  4.120 1.960 5.915 2.285 ;
        RECT  4.595 1.960 5.915 2.300 ;
        RECT  5.685 1.960 5.915 2.350 ;
        RECT  2.850 2.550 4.885 2.845 ;
        RECT  4.595 1.960 4.885 2.845 ;
        RECT  1.555 2.705 3.080 2.935 ;
        RECT  1.555 2.705 1.785 3.090 ;
        RECT  1.865 0.705 4.810 0.935 ;
        RECT  1.865 0.705 2.165 1.390 ;
        RECT  1.490 1.120 2.165 1.390 ;
        RECT  4.580 0.705 4.810 1.730 ;
        RECT  4.580 1.500 8.995 1.730 ;
        RECT  6.750 1.500 8.995 1.870 ;
        RECT  6.750 1.500 7.045 2.850 ;
        RECT  5.450 2.580 7.045 2.850 ;
        RECT  2.390 3.165 2.745 3.510 ;
        RECT  3.310 3.110 5.680 3.340 ;
        RECT  5.450 2.580 5.680 3.340 ;
        RECT  2.390 3.230 3.535 3.510 ;
    END
END BUFT_X16_18_SVT_WB

MACRO BUFT_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN BUFT_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.527  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.885 1.790 4.410 2.130 ;
        RECT  3.885 1.790 4.150 2.395 ;
        END
    END A
    PIN OE
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.915 0.905 2.265 ;
        RECT  0.140 1.730 0.460 2.265 ;
        END
    END OE
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.240  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.435 2.460 8.840 3.290 ;
        RECT  8.485 0.580 8.840 3.290 ;
        RECT  5.645 1.045 8.840 1.300 ;
        RECT  8.405 0.580 8.840 1.300 ;
        RECT  5.715 2.460 8.840 2.775 ;
        RECT  6.985 2.460 7.345 3.290 ;
        RECT  6.960 0.585 7.345 1.300 ;
        RECT  5.715 2.460 7.345 2.780 ;
        RECT  5.645 0.570 6.020 1.300 ;
        RECT  5.715 2.460 5.945 3.290 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  7.700 3.100 8.040 4.100 ;
        RECT  0.825 3.490 1.190 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  7.700 -0.180 8.040 0.760 ;
        RECT  0.655 -0.180 0.995 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.250 0.410 1.605 0.705 ;
        RECT  0.235 0.590 1.365 0.820 ;
        RECT  0.235 0.590 0.465 1.145 ;
        RECT  2.275 2.140 2.560 2.420 ;
        RECT  1.135 2.190 2.560 2.420 ;
        RECT  1.165 0.505 1.365 2.825 ;
        RECT  1.135 0.590 1.365 2.825 ;
        RECT  0.330 2.595 1.365 2.825 ;
        RECT  0.330 2.595 0.560 3.035 ;
        RECT  2.315 1.220 2.655 1.560 ;
        RECT  2.315 1.330 4.870 1.560 ;
        RECT  3.130 2.600 3.360 2.880 ;
        RECT  4.450 2.600 4.870 2.880 ;
        RECT  4.640 1.330 4.870 2.880 ;
        RECT  1.595 2.650 4.870 2.880 ;
        RECT  1.595 2.650 1.935 2.980 ;
        RECT  3.130 0.710 3.360 1.100 ;
        RECT  4.450 0.710 4.680 1.100 ;
        RECT  1.865 0.760 5.330 0.990 ;
        RECT  3.130 0.760 5.330 1.100 ;
        RECT  1.595 0.935 2.090 1.165 ;
        RECT  1.595 0.935 1.880 1.215 ;
        RECT  5.100 1.550 7.890 1.850 ;
        RECT  5.100 0.760 5.330 3.340 ;
        RECT  2.315 3.110 5.330 3.340 ;
        RECT  2.315 3.110 2.600 3.390 ;
    END
END BUFT_X12_18_SVT_WB

MACRO AOI33_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI33_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.660 3.220 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.210 3.800 1.960 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.030 1.565 4.440 2.150 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.095 1.795 2.440 2.150 ;
        RECT  2.095 0.700 2.325 2.150 ;
        RECT  1.770 0.700 2.325 1.085 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.680 1.760 2.150 ;
        RECT  1.250 1.110 1.480 2.150 ;
        RECT  1.030 1.110 1.480 1.450 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.555 1.680 1.020 2.150 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.740 0.535 7.175 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.980 3.515 6.320 4.100 ;
        RECT  1.620 3.070 1.960 4.100 ;
        RECT  0.180 2.440 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.980 -0.180 6.320 0.875 ;
        RECT  4.450 -0.180 4.790 0.405 ;
        RECT  0.460 -0.180 0.800 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.380 2.680 2.720 ;
        RECT  2.340 2.380 2.680 3.190 ;
        RECT  2.340 2.895 4.120 3.190 ;
        RECT  2.560 0.635 4.900 0.975 ;
        RECT  4.670 1.860 5.800 2.180 ;
        RECT  3.060 2.380 4.900 2.665 ;
        RECT  4.670 0.635 4.900 3.410 ;
        RECT  4.500 2.380 4.900 3.410 ;
        RECT  5.220 0.535 5.560 1.485 ;
        RECT  5.220 1.255 6.510 1.485 ;
        RECT  6.280 1.255 6.510 2.750 ;
        RECT  5.220 2.410 6.510 2.750 ;
        RECT  5.220 2.410 5.560 3.385 ;
    END
END AOI33_X4_18_SVT_WB

MACRO AOI33_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI33_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.730 1.660 3.220 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.210 3.800 1.590 ;
        RECT  3.450 1.210 3.725 1.960 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.030 1.565 4.440 2.150 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.095 1.795 2.440 2.150 ;
        RECT  2.095 0.700 2.325 2.150 ;
        RECT  1.770 0.700 2.325 1.085 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.250 1.680 1.760 2.150 ;
        RECT  1.250 1.110 1.480 2.150 ;
        RECT  1.030 1.110 1.480 1.450 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.555 1.680 1.020 2.150 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.940  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.500 2.380 4.900 3.410 ;
        RECT  4.670 0.635 4.900 3.410 ;
        RECT  2.560 0.635 4.900 0.975 ;
        RECT  3.060 2.380 4.900 2.665 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  1.620 3.070 1.960 4.100 ;
        RECT  0.180 2.440 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.450 -0.180 4.790 0.405 ;
        RECT  0.460 -0.180 0.800 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.380 2.680 2.720 ;
        RECT  2.340 2.380 2.680 3.190 ;
        RECT  2.340 2.895 4.120 3.190 ;
    END
END AOI33_X2_18_SVT_WB

MACRO AOI33_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI33_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.375 1.090 2.755 1.625 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.820 3.500 2.265 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.090 4.100 1.590 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.730 1.770 2.180 2.220 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.090 1.660 1.540 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.575 1.690 1.030 2.135 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.870  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 2.535 4.900 2.875 ;
        RECT  4.620 0.615 4.900 2.875 ;
        RECT  2.220 0.615 4.900 0.860 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  1.500 2.450 1.840 4.100 ;
        RECT  0.180 3.110 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.380 -0.180 4.720 0.385 ;
        RECT  0.310 -0.180 0.650 0.930 ;
        END
    END VSS
END AOI33_X1_18_SVT_WB

MACRO AOI33_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI33_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 2.380 2.885 2.720 ;
        RECT  2.545 1.800 2.885 2.720 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.290 1.240 3.830 1.670 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.790 1.900 4.345 2.355 ;
        RECT  4.060 1.715 4.345 2.355 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.815 1.660 2.215 2.165 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.405 0.700 1.745 1.430 ;
        RECT  1.200 0.700 1.745 0.980 ;
        END
    END B1
    PIN B2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.600 1.160 1.050 1.610 ;
        END
    END B2
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.699  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.115 3.050 4.900 3.390 ;
        RECT  4.620 0.625 4.900 3.390 ;
        RECT  2.355 0.625 4.900 0.930 ;
        RECT  3.115 2.380 3.415 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  1.635 2.395 1.975 4.100 ;
        RECT  0.195 3.050 0.535 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.475 -0.180 4.815 0.390 ;
        RECT  0.445 -0.180 0.785 0.930 ;
        END
    END VSS
END AOI33_X0_18_SVT_WB

MACRO AOI32_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI32_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.985 1.820 2.710 2.275 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.170 1.230 3.550 2.100 ;
        RECT  1.260 1.230 3.550 1.590 ;
        RECT  1.260 1.230 1.600 1.960 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.520 2.505 4.330 2.825 ;
        RECT  3.990 1.860 4.330 2.825 ;
        RECT  0.520 1.720 0.860 2.825 ;
        RECT  0.130 1.720 0.860 2.280 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.865 1.175 6.245 1.905 ;
        RECT  5.595 1.175 6.245 1.580 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.020 2.135 7.215 2.365 ;
        RECT  6.745 1.790 7.215 2.365 ;
        RECT  5.020 1.860 5.305 2.365 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.460  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.560 2.595 6.935 2.825 ;
        RECT  2.220 0.635 6.215 0.865 ;
        RECT  5.875 0.470 6.215 0.865 ;
        RECT  4.560 0.635 4.790 2.825 ;
        RECT  2.220 0.635 4.790 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  2.255 3.550 2.605 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  7.025 -0.180 7.365 1.280 ;
        RECT  4.325 -0.180 4.665 0.405 ;
        RECT  0.180 -0.180 0.480 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  7.315 2.595 7.655 3.320 ;
        RECT  0.180 3.055 7.655 3.320 ;
    END
END AOI32_X4_18_SVT_WB

MACRO AOI32_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI32_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.860 2.185 2.710 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.260 1.590 1.965 ;
        RECT  1.010 1.260 1.590 1.540 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.470 1.770 0.980 2.170 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.875 1.260 3.390 1.590 ;
        RECT  2.875 1.260 3.160 1.960 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 1.820 4.020 2.100 ;
        RECT  3.670 1.695 4.020 2.100 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.415 2.380 3.530 2.720 ;
        RECT  2.380 0.550 2.770 1.055 ;
        RECT  2.415 0.550 2.645 2.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  1.710 3.515 2.050 4.100 ;
        RECT  0.230 2.475 0.570 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.915 -0.180 4.255 1.440 ;
        RECT  0.230 -0.180 0.570 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.950 2.475 1.290 3.285 ;
        RECT  3.910 2.495 4.250 3.285 ;
        RECT  0.950 3.015 4.250 3.285 ;
    END
END AOI32_X2_18_SVT_WB

MACRO AOI32_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI32_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.720 1.770 2.170 2.200 ;
        RECT  1.720 1.670 2.050 2.200 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.700 1.610 1.450 ;
        RECT  1.150 0.700 1.610 1.040 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.395 1.260 1.040 1.590 ;
        RECT  0.395 1.105 0.920 1.590 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 1.125 2.770 1.540 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.460 0.650 3.780 1.530 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.830 2.330 3.230 2.720 ;
        RECT  3.000 0.585 3.230 2.720 ;
        RECT  2.115 0.585 3.230 0.890 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.500 2.430 1.840 4.100 ;
        RECT  0.180 3.110 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.395 -0.180 3.740 0.355 ;
        RECT  0.180 -0.180 0.520 0.875 ;
        END
    END VSS
END AOI32_X1_18_SVT_WB

MACRO AOI32_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI32_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.610 1.735 2.125 2.205 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.270 0.700 1.610 1.480 ;
        RECT  1.145 0.700 1.610 1.015 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.410 1.180 0.980 1.665 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.355 1.210 2.710 1.745 ;
        RECT  2.020 1.210 2.710 1.505 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.455 1.055 3.805 1.715 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.830 2.380 3.220 2.720 ;
        RECT  2.940 0.625 3.220 2.720 ;
        RECT  2.180 0.625 3.220 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.510 2.435 1.850 4.100 ;
        RECT  0.180 3.050 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.400 -0.180 3.740 0.370 ;
        RECT  0.180 -0.180 0.530 0.925 ;
        END
    END VSS
END AOI32_X0_18_SVT_WB

MACRO AOI31_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI31_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.770 2.950 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 2.380 3.520 2.770 ;
        RECT  3.180 1.860 3.520 2.770 ;
        RECT  1.810 1.840 2.040 2.770 ;
        RECT  1.190 1.840 2.040 2.180 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.731  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.795 1.860 4.135 2.155 ;
        RECT  3.795 1.260 4.055 2.155 ;
        RECT  0.300 1.260 4.055 1.540 ;
        RECT  0.300 1.260 0.640 1.960 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.535 1.210 5.125 1.680 ;
        RECT  4.535 1.210 4.765 1.960 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.761  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.835 2.515 5.775 2.830 ;
        RECT  5.495 0.640 5.775 2.830 ;
        RECT  2.085 0.640 5.775 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  0.720 3.505 1.085 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  5.490 -0.180 5.835 0.360 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.440 1.580 2.685 ;
        RECT  1.350 2.440 1.580 3.340 ;
        RECT  4.140 2.430 4.480 3.340 ;
        RECT  1.350 3.075 5.925 3.340 ;
    END
END AOI31_X4_18_SVT_WB

MACRO AOI31_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI31_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.960 1.200 2.305 1.960 ;
        RECT  1.820 1.200 2.305 1.610 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.290 1.260 1.590 1.960 ;
        RECT  1.140 1.260 1.590 1.600 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.570 1.820 1.030 2.100 ;
        RECT  0.570 1.570 0.910 2.100 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.320 3.060 2.660 ;
        RECT  2.760 1.840 3.060 2.660 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.119  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.640 3.630 3.375 ;
        RECT  2.570 0.640 3.630 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.810 3.510 2.150 4.100 ;
        RECT  0.330 2.565 0.670 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.330 -0.180 3.670 0.405 ;
        RECT  0.330 -0.180 0.670 1.340 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.050 3.030 2.910 3.265 ;
    END
END AOI31_X2_18_SVT_WB

MACRO AOI31_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI31_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.760 0.690 2.045 1.880 ;
        RECT  1.210 0.690 2.045 1.030 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.260 1.430 1.880 ;
        RECT  0.650 1.260 1.430 1.600 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.125 2.330 0.800 2.710 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.580 2.780 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.581  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 2.890 3.240 3.295 ;
        RECT  3.010 0.995 3.240 3.295 ;
        RECT  2.325 0.995 3.240 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.520 2.535 1.860 4.100 ;
        RECT  0.180 2.955 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.635 -0.180 2.975 0.460 ;
        RECT  0.220 -0.180 0.560 0.460 ;
        END
    END VSS
END AOI31_X1_18_SVT_WB

MACRO AOI31_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI31_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.710 1.770 2.100 2.265 ;
        RECT  1.710 1.720 2.050 2.265 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 0.700 1.600 1.500 ;
        RECT  1.135 0.700 1.600 1.005 ;
        END
    END A1
    PIN A2
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.180 0.980 1.610 ;
        END
    END A2
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.250 1.210 2.785 1.590 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 2.270 3.245 2.780 ;
        RECT  3.015 0.640 3.245 2.780 ;
        RECT  2.280 0.640 3.245 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.500 2.495 1.840 4.100 ;
        RECT  0.180 3.110 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.170 -0.180 0.535 0.920 ;
        END
    END VSS
END AOI31_X0_18_SVT_WB

MACRO AOI22_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI22_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.560 1.210 4.900 1.910 ;
        RECT  4.365 1.210 4.900 1.550 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.820 5.975 2.200 ;
        RECT  4.020 2.140 5.470 2.370 ;
        RECT  3.745 1.860 4.250 2.200 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.605 2.150 2.100 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.800 2.330 3.055 2.560 ;
        RECT  2.715 1.860 3.055 2.560 ;
        RECT  0.800 1.820 1.030 2.560 ;
        RECT  0.650 1.820 1.030 2.205 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.780 2.600 5.860 2.915 ;
        RECT  1.720 0.640 5.020 0.980 ;
        RECT  3.285 2.575 3.895 2.815 ;
        RECT  3.285 0.640 3.515 2.815 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.720 4.100 ;
        RECT  2.480 3.515 2.820 4.100 ;
        RECT  0.960 3.515 1.300 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.720 0.180 ;
        RECT  5.830 -0.180 6.170 1.280 ;
        RECT  3.160 -0.180 3.500 0.405 ;
        RECT  0.570 -0.180 0.910 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 2.520 0.535 3.285 ;
        RECT  0.200 3.045 3.580 3.285 ;
        RECT  6.120 2.385 6.460 3.440 ;
        RECT  3.240 3.155 6.460 3.440 ;
    END
END AOI22_X4_18_SVT_WB

MACRO AOI22_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI22_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.255 0.700 2.770 1.040 ;
        RECT  2.255 0.700 2.540 2.145 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.260 3.270 1.960 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.615 2.300 1.515 2.710 ;
        RECT  1.220 1.840 1.515 2.710 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.560 0.890 1.960 ;
        RECT  0.140 1.145 0.540 1.960 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.750 2.380 2.760 2.720 ;
        RECT  1.750 0.625 2.025 2.720 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.940 3.565 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.140 -0.180 3.480 0.810 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.140 2.475 3.480 3.325 ;
        RECT  0.180 3.015 3.480 3.325 ;
    END
END AOI22_X2_18_SVT_WB

MACRO AOI22_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI22_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.400 1.135 2.160 1.555 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 0.650 3.220 1.545 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.115 1.805 1.620 2.410 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.435 1.150 1.030 1.540 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.594  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.295 2.735 2.945 ;
        RECT  2.390 2.290 2.735 2.945 ;
        RECT  2.390 0.590 2.620 2.945 ;
        RECT  1.685 0.590 2.620 0.820 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.790 3.515 1.140 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.235 -0.180 0.465 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.235 2.660 1.895 2.890 ;
    END
END AOI22_X1_18_SVT_WB

MACRO AOI22_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI22_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.400 1.135 2.160 1.555 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.860 0.650 3.220 1.545 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.115 1.805 1.620 2.290 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.435 1.150 1.030 1.540 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.454  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 2.350 2.735 2.825 ;
        RECT  2.390 2.345 2.735 2.825 ;
        RECT  2.390 0.590 2.620 2.825 ;
        RECT  1.685 0.590 2.620 0.820 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.790 3.515 1.140 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.235 -0.180 0.465 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.235 2.540 1.895 2.770 ;
    END
END AOI22_X0_18_SVT_WB

MACRO AOI222_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI222_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.450 1.820 9.360 2.180 ;
        RECT  7.420 2.180 8.790 2.410 ;
        RECT  6.820 1.840 7.650 2.180 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.880 1.250 8.450 1.590 ;
        RECT  7.880 1.250 8.220 1.950 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.010 2.135 6.440 2.365 ;
        RECT  6.140 1.830 6.440 2.365 ;
        RECT  4.010 1.820 4.390 2.365 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.130 1.260 5.510 1.905 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 2.135 3.140 2.365 ;
        RECT  2.855 1.860 3.140 2.365 ;
        RECT  0.650 1.820 1.030 2.365 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.210 2.200 1.905 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.119  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.330 2.640 9.940 2.880 ;
        RECT  9.600 1.360 9.940 2.880 ;
        RECT  9.240 1.360 9.940 1.590 ;
        RECT  9.240 0.610 9.580 1.590 ;
        RECT  0.455 0.610 9.580 0.865 ;
        RECT  6.635 0.610 6.985 1.390 ;
        RECT  0.455 0.610 0.820 1.400 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  3.060 3.110 3.400 4.100 ;
        RECT  1.620 3.065 1.960 4.100 ;
        RECT  0.180 2.595 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  7.945 -0.180 8.310 0.380 ;
        RECT  5.080 -0.180 5.460 0.350 ;
        RECT  1.660 -0.180 2.000 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.595 6.260 2.835 ;
        RECT  2.340 2.595 6.260 2.880 ;
        RECT  0.900 2.595 1.240 3.405 ;
        RECT  2.340 2.595 2.680 3.405 ;
        RECT  6.625 2.620 6.990 3.450 ;
        RECT  3.760 3.110 9.860 3.450 ;
    END
END AOI222_X4_18_SVT_WB

MACRO AOI222_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI222_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.875 1.685 5.485 2.155 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.805 1.260 4.100 1.960 ;
        RECT  3.385 1.260 4.100 1.540 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.115 1.710 2.700 2.150 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.930 1.850 3.490 2.245 ;
        RECT  2.930 1.735 3.260 2.245 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.380 1.260 1.720 1.960 ;
        RECT  1.120 1.260 1.720 1.540 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.770 1.020 2.240 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.259  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.625 0.630 5.395 0.905 ;
        RECT  4.330 0.630 4.990 1.030 ;
        RECT  4.330 0.630 4.645 2.815 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  0.140 3.055 0.555 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  3.400 -0.180 3.740 0.400 ;
        RECT  0.460 -0.180 0.800 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.475 3.220 2.815 ;
        RECT  0.900 2.475 1.240 3.385 ;
        RECT  5.040 2.385 5.380 3.385 ;
        RECT  2.160 3.045 5.380 3.385 ;
    END
END AOI222_X2_18_SVT_WB

MACRO AOI222_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI222_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.550 1.630 4.925 2.430 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.020 1.230 3.835 1.570 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.770 2.475 2.260 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.790 1.800 3.380 2.205 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.695 1.590 2.205 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.545 0.800 2.210 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.919  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.480 0.590 4.820 1.000 ;
        RECT  3.975 2.415 4.320 2.775 ;
        RECT  4.090 0.590 4.320 2.775 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  0.140 3.405 1.645 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.055 -0.180 3.425 0.360 ;
        RECT  0.220 -0.180 0.530 0.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.750 2.490 2.940 2.775 ;
    END
END AOI222_X1_18_SVT_WB

MACRO AOI222_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI222_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.475 1.755 4.925 2.270 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.230 1.145 3.665 1.540 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 1.820 2.475 2.260 ;
        RECT  2.060 1.770 2.475 2.260 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.790 1.800 3.675 2.205 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.140 1.745 1.590 ;
        END
    END C0
    PIN C1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.160  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.580 1.090 0.995 1.605 ;
        END
    END C1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.714  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.480 0.590 4.820 0.840 ;
        RECT  3.975 0.590 4.385 1.085 ;
        RECT  3.975 0.590 4.205 2.775 ;
        RECT  1.480 0.590 4.385 0.850 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  0.140 3.405 1.645 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.055 -0.180 3.425 0.360 ;
        RECT  0.350 -0.180 0.660 0.430 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.750 2.490 2.940 2.775 ;
    END
END AOI222_X0_18_SVT_WB

MACRO AOI221_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI221_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.175 2.135 7.695 2.365 ;
        RECT  7.385 1.855 7.695 2.365 ;
        RECT  5.175 1.735 5.655 2.365 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.040 1.250 6.670 1.905 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.860 2.980 2.150 ;
        RECT  0.435 2.135 2.685 2.365 ;
        RECT  0.435 1.770 1.050 2.365 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.660 1.260 2.225 1.570 ;
        RECT  1.660 1.260 2.050 1.905 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.340 1.700 4.000 2.115 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 4.213  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.695 2.595 8.265 2.880 ;
        RECT  7.925 1.090 8.265 2.880 ;
        RECT  7.585 0.675 8.010 1.440 ;
        RECT  0.175 0.675 8.010 1.015 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  2.840 3.060 3.185 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  6.355 -0.180 6.705 0.360 ;
        RECT  4.155 -0.180 4.515 0.360 ;
        RECT  1.525 -0.180 1.865 0.350 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.000 2.400 4.615 2.670 ;
        RECT  0.715 2.595 3.295 2.830 ;
        RECT  0.715 2.595 2.465 2.880 ;
        RECT  0.715 2.595 1.095 3.450 ;
        RECT  2.050 2.595 2.465 3.450 ;
        RECT  3.550 3.110 8.225 3.450 ;
    END
END AOI221_X4_18_SVT_WB

MACRO AOI221_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI221_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.750 2.330 4.340 2.710 ;
        RECT  3.750 1.860 4.090 2.710 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.620 1.840 3.060 2.180 ;
        RECT  2.330 2.320 2.850 2.660 ;
        RECT  2.620 1.840 2.850 2.660 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.770 1.720 2.230 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.260 1.135 1.565 ;
        RECT  0.650 1.260 1.000 1.960 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.050 1.260 2.390 1.960 ;
        RECT  1.770 1.260 2.390 1.540 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.692  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.290 0.640 3.970 0.980 ;
        RECT  3.080 2.410 3.520 2.750 ;
        RECT  3.290 0.640 3.520 2.750 ;
        RECT  1.620 0.640 3.970 0.875 ;
        RECT  1.620 0.535 1.960 0.875 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  0.900 3.100 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  2.380 -0.180 2.720 0.405 ;
        RECT  0.470 -0.180 0.810 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.160 2.460 1.980 2.745 ;
        RECT  0.160 2.460 0.520 3.220 ;
        RECT  1.620 2.460 1.980 3.220 ;
        RECT  2.340 3.100 4.120 3.440 ;
    END
END AOI221_X2_18_SVT_WB

MACRO AOI221_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI221_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.860 3.805 2.810 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.590 2.725 2.150 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.770 1.390 2.255 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.590 1.190 1.190 1.540 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.685 1.210 2.115 1.730 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.846  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.675 3.730 0.995 ;
        RECT  2.720 2.380 3.185 2.720 ;
        RECT  2.955 0.675 3.185 2.720 ;
        RECT  1.520 0.675 3.730 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.800 2.485 1.140 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.350 -0.180 0.690 0.930 ;
        END
    END VSS
END AOI221_X1_18_SVT_WB

MACRO AOI221_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI221_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.660 3.805 2.250 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.350 1.660 2.725 2.200 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.155 1.145 1.550 1.675 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.120 1.615 0.770 2.000 ;
        RECT  0.120 1.615 0.430 2.240 ;
        END
    END B1
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.780 1.145 2.195 1.485 ;
        RECT  1.780 1.145 2.115 1.675 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.655  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.955 0.590 3.745 0.930 ;
        RECT  2.810 2.880 3.375 3.260 ;
        RECT  2.810 2.425 3.185 3.260 ;
        RECT  2.955 0.590 3.185 3.260 ;
        RECT  1.370 0.590 3.745 0.915 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.890 2.380 1.230 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  0.220 -0.180 0.520 0.930 ;
        END
    END VSS
END AOI221_X0_18_SVT_WB

MACRO AOI21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.523  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.740 2.145 4.390 2.375 ;
        RECT  3.970 1.790 4.390 2.375 ;
        RECT  1.740 1.915 2.080 2.375 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.523  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.620 1.860 5.605 2.200 ;
        RECT  4.620 1.000 4.935 2.200 ;
        RECT  1.235 1.000 4.935 1.230 ;
        RECT  2.580 1.000 2.920 1.915 ;
        RECT  0.575 1.620 1.510 1.960 ;
        RECT  1.235 1.000 1.510 1.960 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.584  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.955 1.690 7.175 2.225 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.510  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.180 2.535 7.960 2.840 ;
        RECT  7.620 0.470 7.960 2.840 ;
        RECT  7.405 0.995 7.960 2.840 ;
        RECT  5.570 0.995 7.960 1.225 ;
        RECT  6.195 0.460 6.510 1.225 ;
        RECT  5.570 0.540 5.800 1.225 ;
        RECT  1.500 0.540 5.800 0.770 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.960 4.100 ;
        RECT  3.570 3.530 3.925 4.100 ;
        RECT  0.740 3.560 1.080 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.960 0.180 ;
        RECT  8.340 -0.180 8.680 1.280 ;
        RECT  6.900 -0.180 7.240 0.755 ;
        RECT  0.350 -0.180 0.690 1.390 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.640 5.810 2.880 ;
        RECT  5.460 2.640 5.810 3.410 ;
        RECT  1.505 2.640 1.840 3.400 ;
        RECT  2.825 2.640 3.160 3.405 ;
        RECT  8.340 2.600 8.680 3.410 ;
        RECT  5.460 3.070 8.680 3.410 ;
    END
END AOI21_X8_18_SVT_WB

MACRO AOI21_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI21_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.860 2.135 4.390 2.365 ;
        RECT  3.650 1.820 4.390 2.365 ;
        RECT  1.860 1.915 2.200 2.365 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.530 1.455 2.870 1.905 ;
        RECT  1.290 1.455 2.870 1.685 ;
        RECT  0.690 1.675 1.630 2.100 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.620 1.730 5.105 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.178  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.740 2.195 7.080 3.190 ;
        RECT  5.335 2.195 7.080 2.425 ;
        RECT  1.615 0.995 6.335 1.225 ;
        RECT  5.995 0.505 6.335 1.225 ;
        RECT  5.730 0.995 6.070 2.425 ;
        RECT  5.335 2.195 5.640 2.720 ;
        RECT  4.290 0.475 4.630 1.225 ;
        RECT  1.615 0.485 1.965 1.225 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.280 4.100 ;
        RECT  3.820 3.515 4.160 4.100 ;
        RECT  2.340 3.065 2.680 4.100 ;
        RECT  0.900 3.065 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.280 0.180 ;
        RECT  6.750 -0.180 7.105 0.875 ;
        RECT  5.275 -0.180 5.615 0.760 ;
        RECT  3.060 -0.180 3.400 0.765 ;
        RECT  0.470 -0.180 0.810 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.595 4.920 2.835 ;
        RECT  4.580 2.595 4.920 3.385 ;
        RECT  3.060 2.595 3.400 3.385 ;
        RECT  6.020 2.655 6.360 3.385 ;
        RECT  4.580 3.045 6.360 3.385 ;
        RECT  0.180 2.595 0.520 3.405 ;
        RECT  1.620 2.595 1.960 3.405 ;
    END
END AOI21_X6_18_SVT_WB

MACRO AOI21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.260 1.720 1.905 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.150 1.820 3.160 2.180 ;
        RECT  0.660 2.135 2.490 2.365 ;
        RECT  0.660 1.860 0.980 2.365 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.445 1.620 3.825 2.155 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.755  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.780 2.385 4.285 2.725 ;
        RECT  4.055 0.700 4.285 2.725 ;
        RECT  1.620 0.700 4.285 0.980 ;
        RECT  1.620 0.470 1.960 0.980 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  2.340 3.110 2.680 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.515 -0.180 4.840 1.390 ;
        RECT  3.020 -0.180 3.360 0.405 ;
        RECT  0.470 -0.180 0.810 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.640 3.375 2.880 ;
        RECT  3.045 2.640 3.375 3.415 ;
        RECT  4.515 2.605 4.840 3.415 ;
        RECT  3.045 3.075 4.840 3.415 ;
        RECT  0.180 2.640 0.520 3.450 ;
        RECT  1.620 2.640 1.960 3.450 ;
    END
END AOI21_X4_18_SVT_WB

MACRO AOI21_X3_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI21_X3_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.210 1.735 1.690 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.690 1.920 2.870 2.150 ;
        RECT  2.530 1.810 2.870 2.150 ;
        RECT  0.690 1.770 1.030 2.150 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.592  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.010 1.805 4.565 2.170 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.312  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.590 0.660 4.135 0.980 ;
        RECT  3.545 2.400 4.120 2.710 ;
        RECT  3.545 0.660 3.780 2.710 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  2.340 2.840 2.660 4.100 ;
        RECT  0.900 2.840 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.510 -0.180 4.865 0.810 ;
        RECT  2.810 -0.180 3.150 0.430 ;
        RECT  0.470 -0.180 0.810 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.380 3.120 2.610 ;
        RECT  1.620 2.380 1.960 2.740 ;
        RECT  2.890 2.380 3.120 3.180 ;
        RECT  2.890 2.840 3.345 3.180 ;
        RECT  0.180 2.380 0.520 3.180 ;
        RECT  4.500 2.840 4.840 3.180 ;
        RECT  2.890 2.940 4.840 3.180 ;
    END
END AOI21_X3_18_SVT_WB

MACRO AOI21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.235 1.770 1.690 2.265 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.260 1.075 1.600 ;
        RECT  0.650 1.260 0.990 1.960 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.210 2.720 1.910 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.119  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.340 2.180 2.680 3.255 ;
        RECT  1.920 2.180 2.680 2.410 ;
        RECT  1.920 0.630 2.150 2.410 ;
        RECT  1.620 0.630 2.150 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.380 -0.180 2.720 0.880 ;
        RECT  0.465 -0.180 0.810 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.640 1.960 2.870 ;
        RECT  0.180 2.640 0.520 3.450 ;
        RECT  1.620 2.640 1.960 3.450 ;
    END
END AOI21_X2_18_SVT_WB

MACRO AOI21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.100 1.220 1.590 1.685 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.170 0.735 1.700 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.212  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.490 1.925 2.105 2.330 ;
        RECT  1.820 1.685 2.105 2.330 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.634  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.335 1.225 2.660 2.920 ;
        RECT  1.830 1.225 2.660 1.455 ;
        RECT  1.830 0.720 2.060 1.455 ;
        RECT  1.560 0.720 2.060 0.950 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.735 3.515 1.090 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.290 -0.180 2.625 0.995 ;
        RECT  0.175 -0.180 0.520 0.940 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.635 1.840 2.865 ;
    END
END AOI21_X1_18_SVT_WB

MACRO AOI21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.020 1.465 1.570 2.245 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.085 0.590 1.780 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.800 1.460 2.150 2.250 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.428  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.250 2.675 2.660 3.275 ;
        RECT  2.430 1.000 2.660 3.275 ;
        RECT  1.530 1.000 2.660 1.230 ;
        RECT  1.530 0.485 1.870 1.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.765 3.500 1.120 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  2.250 -0.180 2.590 0.770 ;
        RECT  0.180 -0.180 0.500 0.825 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.210 2.670 1.870 3.015 ;
    END
END AOI21_X0_18_SVT_WB

MACRO AOI211_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI211_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.240 1.210 1.585 1.995 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.275 2.380 2.695 2.660 ;
        RECT  2.410 1.860 2.695 2.660 ;
        RECT  0.275 1.840 0.595 2.660 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.840 2.135 5.560 2.660 ;
        RECT  5.220 1.860 5.560 2.660 ;
        RECT  3.385 2.135 5.560 2.365 ;
        RECT  3.385 1.860 3.670 2.365 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.370 1.260 5.010 1.560 ;
        RECT  4.370 1.260 4.750 1.905 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.409  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.500 0.635 5.350 0.980 ;
        RECT  2.925 2.595 4.595 2.825 ;
        RECT  2.925 0.635 3.155 2.825 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  2.260 3.560 2.600 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  2.730 -0.180 3.070 0.405 ;
        RECT  0.180 -0.180 0.500 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.170 3.055 5.780 3.330 ;
    END
END AOI211_X4_18_SVT_WB

MACRO AOI211_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI211_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.620 1.590 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.336  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.135 1.715 0.740 2.245 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.380 2.150 2.660 ;
        RECT  1.820 1.860 2.050 2.660 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.620 2.765 2.100 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.623  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.855 2.380 3.225 3.190 ;
        RECT  2.995 0.470 3.225 3.190 ;
        RECT  1.385 0.700 3.225 1.280 ;
        RECT  2.650 0.470 3.225 1.280 ;
        RECT  1.385 0.470 1.615 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.820 3.515 1.050 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.175 -0.180 0.520 1.280 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.760 0.520 3.120 ;
        RECT  0.180 2.890 1.865 3.120 ;
    END
END AOI211_X2_18_SVT_WB

MACRO AOI211_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI211_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.110 1.590 1.920 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.145 0.980 1.955 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 2.335 2.280 2.760 ;
        RECT  1.820 1.950 2.115 2.760 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.345 1.110 2.785 1.920 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.811  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.740 2.890 3.245 3.295 ;
        RECT  3.015 0.540 3.245 3.295 ;
        RECT  1.400 0.540 3.245 0.880 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.360 3.460 1.170 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.200 -0.180 0.560 0.875 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.250 2.520 0.590 3.220 ;
        RECT  0.250 2.990 1.930 3.220 ;
        RECT  1.590 2.990 1.930 3.330 ;
    END
END AOI211_X1_18_SVT_WB

MACRO AOI211_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AOI211_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.105 1.665 1.865 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.490 1.350 0.980 2.160 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.755 2.380 2.220 2.820 ;
        END
    END B0
    PIN C0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.310 1.105 2.690 1.865 ;
        END
    END C0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.630  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 3.050 3.220 3.390 ;
        RECT  2.920 0.535 3.220 3.390 ;
        RECT  1.400 0.535 3.220 0.875 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.475 3.510 1.270 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.200 -0.180 0.565 0.860 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.240 2.390 0.580 3.280 ;
        RECT  0.240 3.050 2.030 3.280 ;
        RECT  1.690 3.050 2.030 3.390 ;
    END
END AOI211_X0_18_SVT_WB

MACRO AO22_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO22_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.570 1.260 4.950 1.905 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.450 2.135 5.660 2.365 ;
        RECT  5.320 1.860 5.660 2.365 ;
        RECT  3.450 1.770 3.780 2.365 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.260 1.720 1.905 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 2.135 3.220 2.365 ;
        RECT  2.720 1.770 3.220 2.365 ;
        RECT  0.660 1.860 0.980 2.365 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.439  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.400 2.640 8.740 3.395 ;
        RECT  6.860 0.940 8.680 1.280 ;
        RECT  8.340 0.525 8.680 1.280 ;
        RECT  7.940 0.940 8.570 2.980 ;
        RECT  7.080 2.640 8.740 2.980 ;
        RECT  7.080 2.640 7.420 3.395 ;
        RECT  6.860 0.525 7.240 1.280 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  0.900 3.110 1.240 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  5.920 -0.180 6.260 0.405 ;
        RECT  3.190 -0.180 3.530 0.405 ;
        RECT  0.180 -0.180 0.520 1.385 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.640 3.280 2.880 ;
        RECT  1.620 2.640 3.280 2.980 ;
        RECT  2.940 2.640 3.280 3.450 ;
        RECT  0.180 2.640 0.520 3.395 ;
        RECT  1.620 2.640 1.960 3.395 ;
        RECT  2.940 3.110 6.160 3.450 ;
        RECT  1.620 0.635 6.630 0.975 ;
        RECT  6.390 0.635 6.630 2.880 ;
        RECT  6.390 1.860 7.655 2.200 ;
        RECT  6.390 1.860 6.730 2.880 ;
        RECT  3.660 2.595 6.730 2.880 ;
    END
END AO22_X8_18_SVT_WB

MACRO AO22_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO22_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.260 1.710 1.690 2.180 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.660 1.555 1.000 2.150 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.320 1.755 2.775 2.200 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.160 1.260 3.500 1.960 ;
        RECT  2.890 1.260 3.500 1.540 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.360 1.220 4.950 1.560 ;
        RECT  4.360 0.470 4.700 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  5.080 2.640 5.420 4.100 ;
        RECT  3.640 3.110 3.980 4.100 ;
        RECT  2.160 3.515 2.500 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  5.080 -0.180 5.420 0.810 ;
        RECT  3.600 -0.180 3.940 0.405 ;
        RECT  0.180 -0.180 0.520 1.325 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.900 2.945 3.320 3.230 ;
        RECT  1.700 0.695 4.130 1.030 ;
        RECT  3.845 0.695 4.130 2.715 ;
        RECT  0.180 2.430 4.130 2.715 ;
        RECT  0.180 2.430 0.520 3.450 ;
    END
END AO22_X4_18_SVT_WB

MACRO AO22_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO22_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.170 0.820 1.455 1.680 ;
        RECT  0.700 0.820 1.455 1.160 ;
        RECT  0.700 0.590 1.040 1.160 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.175  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.620 0.840 1.850 ;
        RECT  0.500 1.390 0.840 1.850 ;
        RECT  0.140 1.620 0.480 2.275 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.145 1.340 2.660 2.150 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.890 1.340 3.225 2.150 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.995 0.535 4.340 3.270 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  2.010 3.515 3.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.200 -0.180 3.540 0.405 ;
        RECT  0.185 -0.180 0.470 1.160 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.570 2.775 2.910 3.235 ;
        RECT  1.310 3.005 2.910 3.235 ;
        RECT  1.310 3.005 1.650 3.490 ;
        RECT  1.685 0.770 3.765 1.110 ;
        RECT  3.480 0.770 3.765 2.200 ;
        RECT  1.685 0.770 1.915 2.720 ;
        RECT  0.740 2.380 1.915 2.720 ;
    END
END AO22_X2_18_SVT_WB

MACRO AO22_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO22_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.245 1.465 1.665 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.480 1.500 1.015 2.150 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.375 1.685 2.685 2.600 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.915 2.140 3.415 2.600 ;
        RECT  2.915 1.690 3.220 2.600 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.000 0.880 4.340 3.115 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  2.060 3.515 3.540 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.190 -0.180 3.545 0.415 ;
        RECT  0.300 -0.180 0.710 1.150 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.620 2.830 2.960 3.230 ;
        RECT  1.020 3.000 2.960 3.230 ;
        RECT  1.020 3.000 1.360 3.460 ;
        RECT  1.895 0.815 3.770 1.045 ;
        RECT  1.895 0.815 2.250 1.215 ;
        RECT  3.480 0.815 3.770 1.745 ;
        RECT  1.895 0.815 2.125 2.610 ;
        RECT  0.800 2.380 2.125 2.610 ;
        RECT  0.800 2.380 1.275 2.720 ;
    END
END AO22_X1_18_SVT_WB

MACRO AO22_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO22_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.205 1.820 2.725 2.210 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.415 1.160 3.780 1.920 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.160 2.435 1.590 ;
        END
    END B0
    PIN B1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.130 1.820 1.590 2.150 ;
        RECT  1.290 1.340 1.590 2.150 ;
        END
    END B1
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.420  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 2.940 1.090 3.450 ;
        RECT  0.115 0.590 0.600 0.880 ;
        RECT  0.115 0.590 0.345 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  1.450 3.470 1.790 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  3.415 -0.180 3.740 0.930 ;
        RECT  1.020 -0.180 1.360 0.355 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.830 0.590 3.185 0.930 ;
        RECT  0.830 0.590 1.060 1.340 ;
        RECT  0.575 1.110 0.890 1.920 ;
        RECT  2.955 0.590 3.185 2.750 ;
        RECT  2.820 2.440 3.185 2.750 ;
        RECT  0.790 2.440 2.310 2.710 ;
        RECT  2.080 2.440 2.310 3.490 ;
        RECT  2.080 3.150 3.475 3.490 ;
    END
END AO22_X0_18_SVT_WB

MACRO AO21_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO21_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.320 1.360 3.605 1.975 ;
        RECT  1.260 1.360 3.605 1.590 ;
        RECT  1.260 1.360 1.790 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.170 1.820 2.980 2.150 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.295 0.410 4.635 1.940 ;
        RECT  0.800 0.410 4.635 0.640 ;
        RECT  0.650 1.820 1.030 2.195 ;
        RECT  0.800 0.410 1.030 2.195 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.095 0.590 7.435 3.330 ;
        RECT  5.575 1.760 7.435 2.100 ;
        RECT  5.575 0.590 5.915 3.330 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.835 2.630 8.215 4.100 ;
        RECT  6.335 2.630 6.675 4.100 ;
        RECT  4.815 2.630 5.155 4.100 ;
        RECT  0.210 2.480 0.550 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.815 -0.180 8.210 1.290 ;
        RECT  6.335 -0.180 6.675 1.290 ;
        RECT  4.865 -0.180 5.155 0.875 ;
        RECT  0.275 -0.180 0.570 1.435 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.970 2.480 1.310 3.235 ;
        RECT  0.970 2.950 4.395 3.235 ;
        RECT  1.260 0.870 4.065 1.130 ;
        RECT  3.835 2.170 5.345 2.400 ;
        RECT  5.035 1.860 5.345 2.400 ;
        RECT  3.835 0.870 4.065 2.720 ;
        RECT  1.690 2.380 4.065 2.720 ;
    END
END AO21_X8_18_SVT_WB

MACRO AO21_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO21_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.140 1.770 1.540 2.305 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.260 1.030 1.550 ;
        RECT  0.420 1.260 0.760 1.960 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.860 1.260 2.200 1.960 ;
        RECT  1.690 1.260 2.200 1.590 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.060 0.535 3.400 3.390 ;
        RECT  2.940 2.330 3.400 2.990 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.780 2.580 4.120 4.100 ;
        RECT  2.340 3.110 2.680 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.780 -0.180 4.120 1.345 ;
        RECT  2.165 -0.180 2.505 0.405 ;
        RECT  0.180 -0.180 0.520 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 2.635 0.520 3.445 ;
        RECT  0.180 3.105 1.960 3.445 ;
        RECT  1.380 0.550 1.720 0.890 ;
        RECT  1.380 0.635 2.830 0.890 ;
        RECT  2.480 0.635 2.830 2.080 ;
        RECT  2.480 0.635 2.710 2.875 ;
        RECT  0.900 2.535 2.710 2.875 ;
    END
END AO21_X4_18_SVT_WB

MACRO AO21_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO21_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.820 1.340 2.200 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.095 0.815 1.435 ;
        RECT  0.140 1.095 0.475 1.665 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.690 1.640 2.100 2.150 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.875 0.470 3.220 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.120 3.110 2.460 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.120 -0.180 2.460 0.755 ;
        RECT  0.250 -0.180 0.590 0.865 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.400 0.575 1.740 1.215 ;
        RECT  1.400 0.985 2.645 1.215 ;
        RECT  2.330 0.985 2.645 2.775 ;
        RECT  0.780 2.435 2.645 2.775 ;
    END
END AO21_X2_18_SVT_WB

MACRO AO21_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO21_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.650 1.810 1.370 2.150 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.115 1.120 0.900 1.480 ;
        RECT  0.115 1.120 0.430 1.605 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.240 2.100 1.580 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.760 2.920 3.220 3.260 ;
        RECT  2.880 0.985 3.220 3.260 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.000 3.515 2.340 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.280 -0.180 2.625 0.425 ;
        RECT  0.330 -0.180 0.670 0.460 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.520 0.660 2.650 0.960 ;
        RECT  2.330 0.660 2.650 2.225 ;
        RECT  1.630 1.885 2.650 2.225 ;
        RECT  1.630 1.885 1.970 2.720 ;
        RECT  0.800 2.380 1.970 2.720 ;
    END
END AO21_X1_18_SVT_WB

MACRO AO21_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AO21_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.040 1.820 1.590 2.100 ;
        RECT  1.040 1.595 1.380 2.100 ;
        END
    END A0
    PIN A1
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.120 0.550 1.615 ;
        END
    END A1
    PIN B0
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.670 1.120 2.100 1.590 ;
        END
    END B0
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 0.540 3.220 3.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  2.120 3.050 2.460 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  0.180 -0.180 0.520 0.890 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.520 0.550 2.610 0.890 ;
        RECT  2.330 0.550 2.610 2.720 ;
        RECT  0.800 2.380 2.610 2.720 ;
    END
END AO21_X0_18_SVT_WB

MACRO ANTENNA_18_SVT_WB
    CLASS CORE ;
    FOREIGN ANTENNA_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN I
        DIRECTION INPUT ;
        ANTENNADIFFAREA 1.915  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.415 2.340 0.695 3.270 ;
        RECT  0.420 0.550 0.695 1.480 ;
        RECT  0.140 1.090 0.435 2.730 ;
        END
    END I
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 1.120 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 1.120 0.180 ;
        END
    END VSS
END ANTENNA_18_SVT_WB

MACRO AND4_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND4_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.115 1.455 3.455 1.905 ;
        RECT  2.320 1.455 3.455 1.685 ;
        RECT  2.320 1.210 2.660 1.685 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.395 2.135 4.950 2.365 ;
        RECT  4.395 1.820 4.950 2.365 ;
        RECT  2.395 1.915 2.735 2.365 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.685 2.595 5.470 2.825 ;
        RECT  5.180 1.850 5.470 2.825 ;
        RECT  1.685 1.860 2.025 2.825 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.895 1.250 6.235 1.970 ;
        RECT  4.605 1.250 6.235 1.590 ;
        RECT  4.605 0.995 4.945 1.590 ;
        RECT  2.890 0.995 4.945 1.225 ;
        RECT  2.890 0.640 3.205 1.225 ;
        RECT  0.895 0.640 3.205 0.980 ;
        RECT  0.895 0.640 1.235 2.145 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.555 2.420 8.895 3.450 ;
        RECT  7.115 1.040 8.895 1.345 ;
        RECT  8.555 0.535 8.895 1.345 ;
        RECT  7.115 2.420 8.895 2.715 ;
        RECT  7.980 1.040 8.400 2.715 ;
        RECT  7.115 2.420 7.455 3.450 ;
        RECT  7.115 0.535 7.455 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 10.080 4.100 ;
        RECT  9.275 2.640 9.615 4.100 ;
        RECT  7.835 2.945 8.175 4.100 ;
        RECT  6.395 2.890 6.735 4.100 ;
        RECT  4.915 3.515 5.255 4.100 ;
        RECT  3.395 3.515 3.735 4.100 ;
        RECT  1.875 3.515 2.215 4.100 ;
        RECT  0.380 2.640 0.720 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 10.080 0.180 ;
        RECT  9.275 -0.180 9.615 1.345 ;
        RECT  7.835 -0.180 8.175 0.810 ;
        RECT  6.355 -0.180 6.695 0.405 ;
        RECT  0.380 -0.180 0.665 0.810 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.435 0.470 5.765 0.765 ;
        RECT  5.425 0.680 6.885 1.020 ;
        RECT  6.620 1.850 7.680 2.190 ;
        RECT  6.620 0.680 6.885 2.660 ;
        RECT  5.700 2.380 6.885 2.660 ;
        RECT  1.115 2.380 1.455 3.285 ;
        RECT  1.115 3.055 6.015 3.285 ;
        RECT  2.635 3.055 2.975 3.385 ;
        RECT  4.155 3.055 4.495 3.385 ;
        RECT  5.700 2.380 6.015 3.385 ;
        RECT  5.675 3.055 6.015 3.385 ;
    END
END AND4_X8_18_SVT_WB

MACRO AND4_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND4_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.770 0.670 2.185 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.150 1.210 1.490 1.960 ;
        RECT  0.650 1.210 1.490 1.540 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.810 1.210 2.380 1.540 ;
        RECT  1.810 1.210 2.150 1.960 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.770 2.905 2.180 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  5.080 2.320 5.420 3.450 ;
        RECT  3.675 1.580 5.420 1.870 ;
        RECT  5.080 0.535 5.420 1.870 ;
        RECT  3.675 2.320 5.420 2.660 ;
        RECT  4.415 1.580 4.995 2.660 ;
        RECT  3.675 2.320 3.980 3.385 ;
        RECT  3.675 0.535 3.980 1.870 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.600 4.100 ;
        RECT  4.360 3.110 4.700 4.100 ;
        RECT  2.880 2.945 3.220 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.600 0.180 ;
        RECT  4.360 -0.180 4.700 1.345 ;
        RECT  2.880 -0.180 3.220 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.240 0.490 0.580 0.880 ;
        RECT  0.240 0.635 3.445 0.880 ;
        RECT  3.160 0.635 3.445 2.715 ;
        RECT  0.800 2.410 3.445 2.715 ;
        RECT  0.800 2.410 1.140 3.315 ;
        RECT  2.120 2.410 2.460 3.385 ;
    END
END AND4_X6_18_SVT_WB

MACRO AND4_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND4_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.390 1.660 1.005 2.245 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.235 1.185 1.575 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.160 2.235 1.960 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.295 2.325 2.985 2.665 ;
        RECT  2.620 1.770 2.985 2.665 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.800 1.700 4.490 2.185 ;
        RECT  3.800 0.535 4.140 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  4.540 2.480 4.855 4.100 ;
        RECT  3.040 3.515 3.380 4.100 ;
        RECT  1.520 3.515 1.860 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  4.520 -0.180 4.860 1.345 ;
        RECT  3.040 -0.180 3.380 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.470 0.520 1.325 ;
        RECT  0.180 0.635 3.570 0.865 ;
        RECT  0.180 0.635 0.525 1.325 ;
        RECT  3.335 0.635 3.570 3.150 ;
        RECT  0.760 2.895 3.570 3.150 ;
        RECT  0.760 2.475 1.100 3.385 ;
    END
END AND4_X4_18_SVT_WB

MACRO AND4_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND4_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.530 1.620 0.980 2.265 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.620 1.575 2.275 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.805 1.620 2.305 1.960 ;
        RECT  1.805 1.620 2.225 2.445 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.695 1.695 3.250 2.430 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.287  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.995 0.470 4.345 3.190 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  0.395 3.515 3.500 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  2.960 -0.180 3.300 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.330 1.050 3.765 1.390 ;
        RECT  3.480 1.050 3.765 3.015 ;
        RECT  1.050 2.675 3.765 3.015 ;
    END
END AND4_X2_18_SVT_WB

MACRO AND4_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND4_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.165 1.100 1.540 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.980 1.770 1.540 2.305 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.160 2.150 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.770 2.705 2.235 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.540 3.780 2.875 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.190 3.460 3.005 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  2.600 -0.180 2.940 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.310 0.645 3.210 0.930 ;
        RECT  2.935 0.645 3.210 2.875 ;
        RECT  0.740 2.535 3.210 2.875 ;
    END
END AND4_X1_18_SVT_WB

MACRO AND4_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND4_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.380 1.620 3.545 1.960 ;
        RECT  2.380 1.210 2.660 1.960 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.530 1.095 4.900 1.960 ;
        RECT  2.890 1.095 4.900 1.390 ;
        RECT  2.890 0.745 3.120 1.390 ;
        RECT  1.865 0.745 3.120 0.980 ;
        RECT  1.865 0.745 2.150 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 2.190 5.540 2.420 ;
        RECT  5.200 1.860 5.540 2.420 ;
        RECT  1.210 1.820 1.590 2.420 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.525 2.650 6.210 2.880 ;
        RECT  5.870 1.860 6.210 2.880 ;
        RECT  0.525 1.770 0.980 2.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  9.935 0.535 10.275 3.385 ;
        RECT  7.055 1.575 10.275 2.115 ;
        RECT  8.495 0.535 8.835 3.385 ;
        RECT  7.055 0.535 7.395 3.385 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 11.200 4.100 ;
        RECT  10.675 2.445 10.975 4.100 ;
        RECT  9.215 2.575 9.555 4.100 ;
        RECT  7.775 2.575 8.115 4.100 ;
        RECT  6.295 3.570 6.635 4.100 ;
        RECT  4.775 3.570 5.115 4.100 ;
        RECT  3.255 3.570 3.595 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 11.200 0.180 ;
        RECT  10.670 -0.180 10.980 1.365 ;
        RECT  9.215 -0.180 9.555 1.345 ;
        RECT  7.775 -0.180 8.115 1.345 ;
        RECT  6.295 -0.180 6.635 0.405 ;
        RECT  0.180 -0.180 0.520 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  3.350 0.470 3.635 0.865 ;
        RECT  3.350 0.635 6.825 0.865 ;
        RECT  6.505 0.635 6.825 3.340 ;
        RECT  0.785 3.110 6.825 3.340 ;
        RECT  0.785 3.110 1.125 3.450 ;
        RECT  2.105 3.110 2.445 3.450 ;
        RECT  4.015 3.110 4.355 3.450 ;
        RECT  5.535 3.110 5.875 3.450 ;
    END
END AND4_X12_18_SVT_WB

MACRO AND4_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND4_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.510 1.165 1.100 1.540 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.980 1.770 1.540 2.305 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.645 1.160 2.150 1.560 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.270 1.770 2.705 2.235 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.440 0.620 3.780 2.875 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.920 4.100 ;
        RECT  0.190 3.460 3.005 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.920 0.180 ;
        RECT  2.600 -0.180 2.940 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.310 0.645 3.210 0.930 ;
        RECT  2.935 0.645 3.210 2.875 ;
        RECT  0.740 2.535 3.210 2.875 ;
    END
END AND4_X0_18_SVT_WB

MACRO AND3_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND3_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.330 1.565 2.710 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.500 1.105 3.825 1.960 ;
        RECT  1.560 1.105 3.825 1.335 ;
        RECT  1.560 1.105 1.900 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.055 1.770 4.700 2.180 ;
        RECT  0.895 2.330 4.285 2.560 ;
        RECT  4.055 1.770 4.285 2.560 ;
        RECT  0.895 1.840 1.180 2.560 ;
        RECT  0.840 1.840 1.180 2.180 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.444  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  7.160 2.420 7.500 3.190 ;
        RECT  5.720 1.095 7.500 1.335 ;
        RECT  7.160 0.470 7.500 1.335 ;
        RECT  6.690 1.095 7.230 2.720 ;
        RECT  5.720 2.420 7.500 2.720 ;
        RECT  5.720 2.420 6.060 3.230 ;
        RECT  5.720 0.470 6.060 1.335 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 8.400 4.100 ;
        RECT  7.880 2.640 8.220 4.100 ;
        RECT  6.440 3.095 6.780 4.100 ;
        RECT  4.930 3.560 5.270 4.100 ;
        RECT  3.360 3.560 3.700 4.100 ;
        RECT  1.840 3.560 2.180 4.100 ;
        RECT  0.360 2.575 0.665 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 8.400 0.180 ;
        RECT  7.880 -0.180 8.220 1.280 ;
        RECT  6.440 -0.180 6.780 0.810 ;
        RECT  4.680 -0.180 5.180 0.360 ;
        RECT  0.360 -0.180 0.645 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.600 0.590 5.490 0.875 ;
        RECT  5.205 1.705 6.090 2.115 ;
        RECT  5.205 0.590 5.490 3.025 ;
        RECT  1.080 2.790 5.490 3.025 ;
    END
END AND3_X8_18_SVT_WB

MACRO AND3_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND3_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.440 1.725 0.980 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.585 1.545 2.190 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.655 2.200 2.190 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  4.520 2.640 4.860 3.450 ;
        RECT  3.080 1.200 4.860 1.445 ;
        RECT  4.520 0.470 4.860 1.445 ;
        RECT  3.080 2.640 4.860 2.875 ;
        RECT  3.935 1.200 4.370 2.875 ;
        RECT  3.080 2.640 3.420 3.450 ;
        RECT  3.080 0.535 3.420 1.445 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 5.040 4.100 ;
        RECT  3.800 3.110 4.140 4.100 ;
        RECT  2.360 3.110 2.700 4.100 ;
        RECT  0.920 3.110 1.260 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 5.040 0.180 ;
        RECT  3.800 -0.180 4.140 0.970 ;
        RECT  2.320 -0.180 2.660 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.200 0.870 2.850 1.210 ;
        RECT  0.200 0.630 0.540 1.440 ;
        RECT  2.565 1.745 3.400 2.065 ;
        RECT  2.565 0.870 2.850 2.760 ;
        RECT  0.200 2.420 2.850 2.760 ;
        RECT  0.200 2.420 0.540 3.230 ;
        RECT  1.640 2.420 1.980 3.230 ;
    END
END AND3_X6_18_SVT_WB

MACRO AND3_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND3_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.700 1.770 1.110 2.265 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.460 1.260 1.800 1.960 ;
        RECT  1.210 1.260 1.800 1.560 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 2.320 2.520 2.660 ;
        RECT  2.180 1.840 2.520 2.660 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.365 1.110 3.780 1.590 ;
        RECT  3.220 2.575 3.595 3.385 ;
        RECT  3.365 0.535 3.595 3.385 ;
        RECT  3.220 0.535 3.595 1.390 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.940 2.575 4.280 4.100 ;
        RECT  2.460 3.515 2.800 4.100 ;
        RECT  0.940 3.515 1.280 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.940 -0.180 4.280 0.920 ;
        RECT  2.460 -0.180 2.800 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.690 2.990 1.030 ;
        RECT  0.180 0.470 0.520 1.440 ;
        RECT  2.760 1.620 3.135 1.960 ;
        RECT  0.180 2.385 0.465 3.230 ;
        RECT  2.760 0.690 2.990 3.230 ;
        RECT  0.180 2.890 2.990 3.230 ;
    END
END AND3_X4_18_SVT_WB

MACRO AND3_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND3_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.535 1.210 1.115 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.145 1.820 1.595 2.520 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.520 1.230 2.150 1.590 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 2.380 3.225 3.190 ;
        RECT  2.945 0.535 3.225 3.190 ;
        RECT  2.840 0.535 3.225 1.440 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.940 3.515 2.430 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.080 -0.180 2.420 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.420 0.690 2.610 0.980 ;
        RECT  2.380 1.835 2.715 2.175 ;
        RECT  2.380 0.690 2.610 3.075 ;
        RECT  0.180 2.775 2.610 3.075 ;
    END
END AND3_X2_18_SVT_WB

MACRO AND3_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND3_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 2.205 0.745 2.545 ;
        RECT  0.140 1.770 0.465 2.545 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.090 1.680 1.540 2.150 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.770 1.700 2.100 2.325 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 2.890 3.220 3.270 ;
        RECT  2.990 1.005 3.220 3.270 ;
        RECT  2.800 1.005 3.220 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.940 3.515 2.425 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.040 -0.180 2.380 0.870 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 1.100 2.570 1.440 ;
        RECT  2.340 2.255 2.760 2.595 ;
        RECT  2.340 1.100 2.570 3.115 ;
        RECT  0.180 2.775 2.570 3.115 ;
    END
END AND3_X1_18_SVT_WB

MACRO AND3_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND3_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.030 1.620 2.850 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.245 1.095 3.585 1.960 ;
        RECT  1.220 1.095 3.585 1.390 ;
        RECT  1.220 1.095 1.560 1.960 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.530 2.350 4.360 2.580 ;
        RECT  4.005 1.840 4.360 2.580 ;
        RECT  0.530 1.725 0.990 2.580 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.627  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  8.180 0.470 8.520 3.230 ;
        RECT  5.300 1.680 8.520 2.110 ;
        RECT  6.740 0.470 7.150 3.230 ;
        RECT  5.300 1.680 7.150 2.115 ;
        RECT  5.300 0.470 5.640 3.230 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 9.520 4.100 ;
        RECT  8.900 2.640 9.240 4.100 ;
        RECT  7.460 2.640 7.800 4.100 ;
        RECT  6.020 2.640 6.360 4.100 ;
        RECT  4.540 3.375 4.880 4.100 ;
        RECT  3.020 3.515 3.360 4.100 ;
        RECT  1.500 3.515 1.840 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 9.520 0.180 ;
        RECT  8.900 -0.180 9.240 1.280 ;
        RECT  7.460 -0.180 7.800 0.810 ;
        RECT  6.020 -0.180 6.360 1.280 ;
        RECT  4.425 -0.180 4.765 0.405 ;
        RECT  0.310 -0.180 0.650 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.260 0.470 2.600 0.865 ;
        RECT  2.260 0.635 5.070 0.865 ;
        RECT  4.760 0.635 5.070 3.145 ;
        RECT  0.740 2.905 5.070 3.145 ;
    END
END AND3_X12_18_SVT_WB

MACRO AND3_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND3_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.295 1.205 1.230 1.545 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.820 1.605 2.335 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.835 1.205 2.150 1.780 ;
        RECT  1.770 1.205 2.150 1.545 ;
        END
    END C
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.840 2.630 3.220 2.970 ;
        RECT  2.990 0.650 3.220 2.970 ;
        RECT  2.840 0.650 3.220 1.030 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  0.960 3.515 2.425 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  2.080 -0.180 2.420 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.650 2.610 0.975 ;
        RECT  2.380 1.675 2.760 2.015 ;
        RECT  2.380 0.650 2.610 2.970 ;
        RECT  0.200 2.630 2.610 2.970 ;
    END
END AND3_X0_18_SVT_WB

MACRO AND2_X8_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND2_X8_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.135 1.620 1.590 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.820 1.920 2.810 2.150 ;
        RECT  2.380 1.640 2.810 2.150 ;
        RECT  0.520 2.330 2.050 2.560 ;
        RECT  1.820 1.920 2.050 2.560 ;
        RECT  0.520 1.840 0.860 2.560 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.376  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.700 2.695 5.360 3.395 ;
        RECT  5.020 0.590 5.360 3.395 ;
        RECT  3.500 1.050 5.360 1.345 ;
        RECT  3.500 0.590 3.840 1.345 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 6.160 4.100 ;
        RECT  2.980 3.110 3.320 4.100 ;
        RECT  1.500 3.515 1.840 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 6.160 0.180 ;
        RECT  4.260 -0.180 4.600 0.820 ;
        RECT  2.740 -0.180 3.080 0.820 ;
        RECT  0.310 -0.180 0.650 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.470 0.590 1.810 1.345 ;
        RECT  1.470 1.050 3.270 1.345 ;
        RECT  3.040 1.860 4.485 2.200 ;
        RECT  3.040 1.050 3.270 2.700 ;
        RECT  2.280 2.470 3.270 2.700 ;
        RECT  2.280 2.470 2.600 3.280 ;
        RECT  0.725 3.045 2.600 3.280 ;
    END
END AND2_X8_18_SVT_WB

MACRO AND2_X6_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND2_X6_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.380 1.820 1.060 2.100 ;
        RECT  0.380 1.665 0.940 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.330 1.260 1.660 2.065 ;
        RECT  1.170 1.260 1.660 1.540 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 2.244  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  3.960 2.150 4.300 3.450 ;
        RECT  2.520 1.250 4.300 1.590 ;
        RECT  3.960 0.470 4.300 1.590 ;
        RECT  2.520 2.150 4.300 2.390 ;
        RECT  3.235 1.250 3.795 2.390 ;
        RECT  2.520 2.150 2.860 3.450 ;
        RECT  2.520 0.535 2.860 1.590 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 4.480 4.100 ;
        RECT  3.240 2.640 3.580 4.100 ;
        RECT  1.800 2.890 2.140 4.100 ;
        RECT  0.360 2.480 0.700 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 4.480 0.180 ;
        RECT  3.240 -0.180 3.580 0.810 ;
        RECT  1.760 -0.180 2.100 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.360 0.490 0.720 1.430 ;
        RECT  0.360 0.690 2.290 1.030 ;
        RECT  0.360 0.690 0.730 1.430 ;
        RECT  1.990 0.690 2.290 2.660 ;
        RECT  1.080 2.330 2.290 2.660 ;
        RECT  1.080 2.330 1.420 3.450 ;
    END
END AND2_X6_18_SVT_WB

MACRO AND2_X4_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND2_X4_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.615 0.570 2.150 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.396  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.110 1.720 1.540 2.190 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.188  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.290 0.470 2.780 3.190 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 3.360 4.100 ;
        RECT  1.520 3.110 1.860 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 3.360 0.180 ;
        RECT  1.480 -0.180 1.820 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.190 0.485 0.515 1.335 ;
        RECT  0.190 0.995 2.060 1.335 ;
        RECT  1.770 0.995 2.060 2.760 ;
        RECT  0.800 2.420 2.060 2.760 ;
        RECT  0.800 2.420 1.140 3.230 ;
    END
END AND2_X4_18_SVT_WB

MACRO AND2_X2_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND2_X2_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.140 1.535 0.760 2.205 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.198  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.195 1.255 1.590 1.795 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 1.056  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.325 0.535 2.660 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.180 3.110 0.520 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.520 -0.180 1.860 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.795 2.095 1.025 ;
        RECT  0.180 0.795 0.520 1.135 ;
        RECT  1.820 0.795 2.095 2.975 ;
        RECT  0.900 2.635 2.095 2.975 ;
        RECT  0.900 2.635 1.240 3.295 ;
    END
END AND2_X2_18_SVT_WB

MACRO AND2_X1_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND2_X1_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.465 1.205 0.980 1.600 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.210 1.205 1.590 1.740 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.528  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.280 0.540 2.660 3.260 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.175 3.510 1.860 4.100 ;
        RECT  1.520 2.920 1.860 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.520 -0.180 1.860 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.645 2.050 0.975 ;
        RECT  1.820 0.645 2.050 2.690 ;
        RECT  0.760 2.455 2.050 2.690 ;
        RECT  0.760 2.455 1.100 3.105 ;
    END
END AND2_X1_18_SVT_WB

MACRO AND2_X12_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND2_X12_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.640 1.620 2.100 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.792  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.850 1.820 2.900 2.180 ;
        RECT  0.610 2.330 2.135 2.560 ;
        RECT  1.850 1.820 2.135 2.560 ;
        RECT  0.610 1.860 0.950 2.560 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 3.564  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  6.640 0.470 6.980 3.450 ;
        RECT  5.200 1.820 6.980 2.220 ;
        RECT  5.200 0.470 5.540 3.450 ;
        RECT  3.760 1.820 6.980 2.205 ;
        RECT  3.760 0.470 4.100 3.450 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 7.840 4.100 ;
        RECT  5.920 2.640 6.260 4.100 ;
        RECT  4.480 2.640 4.820 4.100 ;
        RECT  3.040 3.110 3.380 4.100 ;
        RECT  1.560 3.570 1.900 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 7.840 0.180 ;
        RECT  5.920 -0.180 6.260 1.280 ;
        RECT  4.480 -0.180 4.820 1.280 ;
        RECT  2.840 -0.180 3.180 0.875 ;
        RECT  0.180 -0.180 0.520 1.440 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  1.600 0.470 1.940 1.410 ;
        RECT  1.600 1.105 3.530 1.410 ;
        RECT  3.230 1.105 3.530 2.750 ;
        RECT  2.365 2.410 3.530 2.750 ;
        RECT  2.365 2.410 2.660 3.340 ;
        RECT  0.800 3.045 2.660 3.340 ;
    END
END AND2_X12_18_SVT_WB

MACRO AND2_X0_18_SVT_WB
    CLASS CORE ;
    FOREIGN AND2_X0_18_SVT_WB 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  0.420 1.210 0.980 1.590 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        ANTENNAMODEL OXIDE1 ;
        ANTENNAGATEAREA 0.151  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  1.180 1.720 1.590 2.355 ;
        END
    END B
    PIN Q
        DIRECTION OUTPUT ;
        ANTENNADIFFAREA 0.403  LAYER M1  ;
        PORT
        LAYER M1 ;
        RECT  2.315 0.540 2.660 3.060 ;
        END
    END Q
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 3.740 2.800 4.100 ;
        RECT  0.195 3.460 1.885 4.100 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER M1 ;
        RECT  0.000 -0.180 2.800 0.180 ;
        RECT  1.520 -0.180 1.860 0.405 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.180 0.540 0.520 0.980 ;
        RECT  0.180 0.750 2.085 0.980 ;
        RECT  1.820 0.750 2.085 3.060 ;
        RECT  0.900 2.720 2.085 3.060 ;
    END
END AND2_X0_18_SVT_WB

END LIBRARY
