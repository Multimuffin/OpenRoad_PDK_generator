/opt/tech/tower/digital/tsl18fs191svt_wb_Rev_2020.03/lib/cdl/tsl18fs191svt_wb.cdl