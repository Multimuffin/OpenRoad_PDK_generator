/opt/tech/tower/digital/tsl18fs190svt_wb_Rev_2022.12/lib/lef/tsl18fs190svt_wb.lef