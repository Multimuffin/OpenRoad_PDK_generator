/opt/tech/tower/digital/tsl18fs190svt_wb_Rev_2022.12/tech/lef/5M1L/tsl180l5.lef