/opt/tech/tower/digital/tsl18fs190svt_Rev_2019.09/tech/lef/6M1L/tsl180l6.lef