*  -------------------------------------- *
* Defining the default unit for both length and area
*.SCALE meter
*  -------------------------------------- *
.option scale=1

.subckt AND2_X0_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q_neg A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q Q_neg VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AND2_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q_neg A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AND2_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD A net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M4 net_000 B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD B Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND2_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND3_X0_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS C net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD B net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD C net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AND3_X1_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_1 B net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS C net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q_neg B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD C Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AND3_X12_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_004 B net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q net_002 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND3_X2_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_1 B net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS C net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M5 Q_neg B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD C Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND3_X4_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_001 A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND3_X6_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND3_X8_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 B net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND4_X0_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_1 B net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_2 C net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS D net_2 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q_neg A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q_neg C VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD D Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q Q_neg VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AND4_X1_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_1 B net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_2 C net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS D net_2 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M5 Q_neg A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q_neg C VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD D Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AND4_X12_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_003 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 A net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_005 B net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_005 C net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS D net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q net_003 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q net_003 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND4_X2_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_1 B net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_2 C net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS D net_2 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q_neg A VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q_neg C VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD D Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND4_X4_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 C net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS D net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD D net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND4_X6_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_0 A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_1 B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_2 C net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS D net_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD B Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q_neg C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD D Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AND4_X8_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_2_1 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_1_1 C net_2_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_1 B net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q_neg A net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_0 A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_1_0 B net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_2_0 C net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS D net_2_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q_neg D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q_neg B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD B Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q_neg C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD D Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt ANTENNA_18_SVT_WB I VDD VSS
*.PININFO I:I VDD:B VSS:B
D0 VSS I DN AREA=0.9156e-12 PJ=3.86e-06
D1 I VDD DP AREA=0.9996e-12 PJ=4.06e-06
.ends

.subckt AO21_X0_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q_neg A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B0 Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q_neg A1 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 A0 Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B0 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AO21_X1_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q_neg A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B0 Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q_neg A1 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 A0 Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B0 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AO21_X2_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q_neg A0 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS B0 Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q_neg A1 net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_1 A0 Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B0 net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AO21_X4_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_001 A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_002 A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AO21_X8_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q_neg B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_0_1 A0 Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A1 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q_neg A0 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B0 Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_1 B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q_neg A0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_1 A1 Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q_neg A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_1 A0 Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AO22_X0_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS net_001 Q VSS N_ISO W=0.455e-06 L=0.18e-06
M1 VSS B1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_001 B0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_001 A0 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS A1 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD net_001 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_003 A0 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_003 A1 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AO22_X1_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q_neg A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_1 B0 Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B1 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_2 A1 Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q_neg A0 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_2 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD B1 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AO22_X2_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_001 A0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 B0 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B1 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_003 A1 net_001 VDD P_ISO W=0.45e-06 L=0.18e-06
M6 net_003 A0 net_001 VDD P_ISO W=0.45e-06 L=0.18e-06
M7 VDD B0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AO22_X4_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_003 A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_001 A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AO22_X8_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A1 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_001 A0 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_001 A0 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A1 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD B1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD B0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_001 A1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_005 A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_001 A0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_001 A1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI211_X0_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q C0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A1 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 A0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_2 B0 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q C0 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI211_X1_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q A0 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS B0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q C0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A1 net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_1 A0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_2 B0 net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q C0 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AOI211_X2_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A0 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q C0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A1 net_1 VDD P_ISO W=0.815e-06 L=0.18e-06
M5 net_1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_2 B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q C0 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI211_X4_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 net_0_0_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A0 net_0_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_0_1 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_0_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q C0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_1 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_2_0_0 B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q C0 net_2_0_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_2_0_1 C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_1 B0 net_2_0_1 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI21_X0_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD A1 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M4 net_1 A0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q B0 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI21_X1_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=0.565e-06 L=0.18e-06
M1 Q A0 net_0 VSS N_ISO W=0.565e-06 L=0.18e-06
M2 VSS B0 Q VSS N_ISO W=0.565e-06 L=0.18e-06
M3 VDD A1 net_1 VDD P_ISO W=0.615e-06 L=0.18e-06
M4 net_1 A0 VDD VDD P_ISO W=0.615e-06 L=0.18e-06
M5 Q B0 net_1 VDD P_ISO W=0.615e-06 L=0.18e-06
.ends

.subckt AOI21_X2_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A0 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 net_1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI21_X3_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0_0_1 A1 VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M1 Q A0 net_0_0_1 VSS N_ISO W=0.785e-06 L=0.18e-06
M2 net_0_0_0 A0 Q VSS N_ISO W=0.785e-06 L=0.18e-06
M3 VSS A1 net_0_0_0 VSS N_ISO W=0.785e-06 L=0.18e-06
M4 Q B0 VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M5 VSS B0 Q VSS N_ISO W=0.785e-06 L=0.18e-06
M6 VDD A1 net_1 VDD P_ISO W=0.86e-06 L=0.18e-06
M7 net_1 A0 VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M8 VDD A0 net_1 VDD P_ISO W=0.86e-06 L=0.18e-06
M9 net_1 A1 VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M10 Q B0 net_1 VDD P_ISO W=0.86e-06 L=0.18e-06
M11 net_1 B0 Q VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt AOI21_X4_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0_1 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A0 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_0 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_1 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_1 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI21_X6_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A0 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_1 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_2 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A0 net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_1 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_1 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI21_X8_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_0_3 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A0 net_0_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_2 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_1 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A0 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_0 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A1 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD A1 net_1 VDD P_ISO W=0.81e-06 L=0.18e-06
M13 net_1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_1 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_1 A0 VDD VDD P_ISO W=0.81e-06 L=0.18e-06
M18 VDD A0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_1 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_1 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 net_1 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI221_X0_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q B0 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS C0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_0 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD B1 net_3 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_3 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_2 C0 net_3 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q A1 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_2 A0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI221_X1_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q B0 net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS C0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_0 A1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q A0 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD B1 net_3 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_3 B0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_2 C0 net_3 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q A1 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_2 A0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AOI221_X2_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q B0 net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A0 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD B1 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_3 B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_2 C0 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q A1 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_2 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI221_X4_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q C0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS A1 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q A0 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_005 C0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_005 C0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q A0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_005 A1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q A1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q A0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI222_X0_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 VSS C1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q C0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q B0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B1 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS A1 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q A0 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VDD C1 net_003 VDD P_ISO W=0.47e-06 L=0.18e-06
M7 VDD C0 net_003 VDD P_ISO W=0.47e-06 L=0.18e-06
M8 net_004 B0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_004 B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 net_004 A1 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M11 net_004 A0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI222_X1_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 VSS C1 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q C0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q B0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B1 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A1 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 Q A0 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VDD C1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD C0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_004 B0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_004 B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_004 A1 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_004 A0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AOI222_X2_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 net_2 C1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q C0 net_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_1 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B1 net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A0 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_4 C1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD C0 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_4 B0 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_3 B1 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q A1 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_3 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI222_X4_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 net_2_0 C0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C1 net_2_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_2_1 C1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q C0 net_2_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_1_0 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B1 net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_1_1 B1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q B0 net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_0 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS A1 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_0_1 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q A0 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_4 C0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C1 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_4 C1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD C0 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_4 B0 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_3 B1 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_4 B1 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_3 B0 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q A0 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_3 A1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q A1 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 net_3 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI22_X0_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q B0 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_0 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS A1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD B1 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_2 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q A0 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_2 A1 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI22_X1_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q B0 net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_0 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS A1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD B1 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_2 B0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q A0 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_2 A1 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AOI22_X2_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q B0 net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD B1 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 net_2 B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q A0 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_2 A1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI22_X4_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1_0 B1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q B0 net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_1_1 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B1 net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_0 A1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A0 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_1 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A1 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD B1 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_2 B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B0 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_2 B1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q A1 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_2 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A0 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_2 A1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI31_X0_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 net_1 A2 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_0 A1 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_2 A2 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD A1 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_2 A0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q B0 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI31_X1_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 net_1 A2 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_0 A1 net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q A0 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_2 A2 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD A1 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_2 A0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q B0 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AOI31_X2_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 net_1 A2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_0 A1 net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A0 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_2 A2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD A1 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_2 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q B0 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI31_X4_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 VSS A2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 A1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A2 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A2 net_004 VDD P_ISO W=0.81e-06 L=0.18e-06
M9 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A2 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_004 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI32_X0_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_2 A2 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_1 A1 net_2 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q A0 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_0 B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS B1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_3 A2 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD A1 net_3 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_3 A0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q B0 net_3 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_3 B1 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI32_X1_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_2 A2 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_1 A1 net_2 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q A0 net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_0 B0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS B1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_3 A2 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD A1 net_3 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_3 A0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B0 net_3 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_3 B1 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AOI32_X2_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_2 A2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_1 A1 net_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A0 net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_3 A2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD A1 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_3 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q B0 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_3 B1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI32_X4_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_2_0 A2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_1_0 A1 net_2_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A0 net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_1_1 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_2_1 A1 net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A2 net_2_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_0 B1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q B0 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_1 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B1 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD A2 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_3 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A0 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_3 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A1 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_3 A2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q B1 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_3 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q B0 net_3 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_3 B1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI33_X0_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 net_3 B2 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_2 B1 net_3 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q B0 net_2 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_0 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_1 A1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS A2 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 net_4 B2 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B1 net_4 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_4 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q A0 net_4 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 net_4 A1 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M11 Q A2 net_4 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt AOI33_X1_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 net_3 B2 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_2 B1 net_3 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q B0 net_2 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_0 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_1 A1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS A2 net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 net_4 B2 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD B1 net_4 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_4 B0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q A0 net_4 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_4 A1 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M11 Q A2 net_4 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt AOI33_X2_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 net_3 B2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_2 B1 net_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q B0 net_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_1 A1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A2 net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_4 B2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B1 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_4 B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A0 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_4 A1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A2 net_4 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt AOI33_X4_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 VSS B2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 A0 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_004 A1 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A2 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_005 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_005 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD B2 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B1 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B0 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_002 A0 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_006 A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_006 A2 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_002 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_005 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_005 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUFT_X1_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE NOE VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_0 NOE VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_1 OE net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS A net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q net_0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD OE NOE VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_1 OE VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_0 NOE net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD A net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q net_1 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt BUFT_X12_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE NOE VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_0 NOE VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M2 net_1 OE net_0 VSS N_ISO W=0.71e-06 L=0.18e-06
M3 net_0 OE net_1 VSS N_ISO W=0.71e-06 L=0.18e-06
M4 VSS A net_0 VSS N_ISO W=0.71e-06 L=0.18e-06
M5 net_0 A VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M6 Q net_0 VSS VSS N_ISO W=0.95e-06 L=0.18e-06
M7 VSS net_0 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M8 Q net_0 VSS VSS N_ISO W=0.95e-06 L=0.18e-06
M9 VSS net_0 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M10 Q net_0 VSS VSS N_ISO W=0.95e-06 L=0.18e-06
M11 VSS net_0 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M12 VDD OE NOE VDD P_ISO W=0.575e-06 L=0.18e-06
M13 net_1 OE VDD VDD P_ISO W=0.78e-06 L=0.18e-06
M14 net_0 NOE net_1 VDD P_ISO W=0.78e-06 L=0.18e-06
M15 net_1 NOE net_0 VDD P_ISO W=0.78e-06 L=0.18e-06
M16 VDD A net_1 VDD P_ISO W=0.755e-06 L=0.18e-06
M17 net_1 A VDD VDD P_ISO W=0.755e-06 L=0.18e-06
M18 Q net_1 VDD VDD P_ISO W=1.05e-06 L=0.18e-06
M19 VDD net_1 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M20 Q net_1 VDD VDD P_ISO W=1.05e-06 L=0.18e-06
M21 VDD net_1 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M22 Q net_1 VDD VDD P_ISO W=1.05e-06 L=0.18e-06
M23 VDD net_1 Q VDD P_ISO W=1.05e-06 L=0.18e-06
.ends

.subckt BUFT_X16_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE net_000 VSS N_ISO W=0.53e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.71e-06 L=0.18e-06
M2 net_001 OE net_002 VSS N_ISO W=0.71e-06 L=0.18e-06
M3 net_001 OE net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_001 VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VSS A net_001 VSS N_ISO W=0.95e-06 L=0.18e-06
M6 VSS A net_001 VSS N_ISO W=0.95e-06 L=0.18e-06
M7 Q net_001 VSS VSS N_ISO W=0.95e-06 L=0.18e-06
M8 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M9 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M10 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M11 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M12 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M13 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M14 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M15 VDD OE net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M16 VDD OE net_002 VDD P_ISO W=0.78e-06 L=0.18e-06
M17 net_002 net_000 net_001 VDD P_ISO W=0.78e-06 L=0.18e-06
M18 net_001 net_000 net_002 VDD P_ISO W=0.86e-06 L=0.18e-06
M19 VDD A net_002 VDD P_ISO W=0.69e-06 L=0.18e-06
M20 VDD A net_002 VDD P_ISO W=0.79e-06 L=0.18e-06
M21 VDD A net_002 VDD P_ISO W=0.79e-06 L=0.18e-06
M22 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M23 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M24 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M25 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M26 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M27 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M28 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M29 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
.ends

.subckt BUFT_X2_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE NOE VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_0 NOE VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_1 OE net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS A net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q net_0 VSS VSS N_ISO W=0.625e-06 L=0.18e-06
M5 VDD OE NOE VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_1 OE VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_0 NOE net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD A net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q net_1 VDD VDD P_ISO W=0.69e-06 L=0.18e-06
.ends

.subckt BUFT_X20_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE NOE VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_0 NOE VSS VSS N_ISO W=0.65e-06 L=0.18e-06
M2 net_1 OE net_0 VSS N_ISO W=0.65e-06 L=0.18e-06
M3 net_0 OE net_1 VSS N_ISO W=0.65e-06 L=0.18e-06
M4 net_1 OE net_0 VSS N_ISO W=0.65e-06 L=0.18e-06
M5 net_0 OE net_1 VSS N_ISO W=0.65e-06 L=0.18e-06
M6 VSS A net_0 VSS N_ISO W=0.65e-06 L=0.18e-06
M7 net_0 A VSS VSS N_ISO W=0.65e-06 L=0.18e-06
M8 VSS A net_0 VSS N_ISO W=0.65e-06 L=0.18e-06
M9 net_0 A VSS VSS N_ISO W=0.65e-06 L=0.18e-06
M10 Q net_0 VSS VSS N_ISO W=0.9e-06 L=0.18e-06
M11 VSS net_0 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M12 Q net_0 VSS VSS N_ISO W=0.9e-06 L=0.18e-06
M13 VSS net_0 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M14 Q net_0 VSS VSS N_ISO W=0.9e-06 L=0.18e-06
M15 VSS net_0 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M16 Q net_0 VSS VSS N_ISO W=0.9e-06 L=0.18e-06
M17 VSS net_0 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M18 Q net_0 VSS VSS N_ISO W=0.9e-06 L=0.18e-06
M19 VSS net_0 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M20 VDD OE NOE VDD P_ISO W=0.575e-06 L=0.18e-06
M21 net_1 OE VDD VDD P_ISO W=0.72e-06 L=0.18e-06
M22 net_0 NOE net_1 VDD P_ISO W=0.72e-06 L=0.18e-06
M23 net_1 NOE net_0 VDD P_ISO W=0.72e-06 L=0.18e-06
M24 net_0 NOE net_1 VDD P_ISO W=0.72e-06 L=0.18e-06
M25 net_1 NOE net_0 VDD P_ISO W=0.72e-06 L=0.18e-06
M26 VDD A net_1 VDD P_ISO W=0.72e-06 L=0.18e-06
M27 net_1 A VDD VDD P_ISO W=0.72e-06 L=0.18e-06
M28 VDD A net_1 VDD P_ISO W=0.72e-06 L=0.18e-06
M29 net_1 A VDD VDD P_ISO W=0.72e-06 L=0.18e-06
M30 Q net_1 VDD VDD P_ISO W=1e-06 L=0.18e-06
M31 VDD net_1 Q VDD P_ISO W=1e-06 L=0.18e-06
M32 Q net_1 VDD VDD P_ISO W=1e-06 L=0.18e-06
M33 VDD net_1 Q VDD P_ISO W=1e-06 L=0.18e-06
M34 Q net_1 VDD VDD P_ISO W=1e-06 L=0.18e-06
M35 VDD net_1 Q VDD P_ISO W=1e-06 L=0.18e-06
M36 Q net_1 VDD VDD P_ISO W=1e-06 L=0.18e-06
M37 VDD net_1 Q VDD P_ISO W=1e-06 L=0.18e-06
M38 Q net_1 VDD VDD P_ISO W=1e-06 L=0.18e-06
M39 VDD net_1 Q VDD P_ISO W=1e-06 L=0.18e-06
.ends

.subckt BUFT_X24_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.65e-06 L=0.18e-06
M2 net_001 OE net_002 VSS N_ISO W=1.055e-06 L=0.18e-06
M3 net_001 OE net_002 VSS N_ISO W=1.055e-06 L=0.18e-06
M4 net_002 OE net_001 VSS N_ISO W=1.055e-06 L=0.18e-06
M5 net_001 OE net_002 VSS N_ISO W=1.055e-06 L=0.18e-06
M6 VSS A net_001 VSS N_ISO W=1.055e-06 L=0.18e-06
M7 VSS A net_001 VSS N_ISO W=1.055e-06 L=0.18e-06
M8 VSS A net_001 VSS N_ISO W=1.055e-06 L=0.18e-06
M9 VSS A net_001 VSS N_ISO W=0.875e-06 L=0.18e-06
M10 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M11 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M12 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M13 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M14 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M15 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M16 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M17 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M18 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M19 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M20 VSS net_001 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M21 VDD OE net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M22 VDD OE net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M23 net_001 net_000 net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M24 net_001 net_000 net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M25 net_001 net_000 net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M26 net_001 net_000 net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M27 VDD A net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M28 VDD A net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M29 VDD A net_002 VDD P_ISO W=0.935e-06 L=0.18e-06
M30 VDD A net_002 VDD P_ISO W=0.72e-06 L=0.18e-06
M31 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M32 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M33 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M34 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M35 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M36 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M37 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M38 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M39 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M40 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
M41 VDD net_002 Q VDD P_ISO W=1e-06 L=0.18e-06
.ends

.subckt BUFT_X3_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 OE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS net_002 Q VSS N_ISO W=0.615e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.615e-06 L=0.18e-06
M6 VDD OE net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD OE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_001 net_000 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_001 A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD net_001 Q VDD P_ISO W=0.7e-06 L=0.18e-06
M11 VDD net_001 Q VDD P_ISO W=0.7e-06 L=0.18e-06
.ends

.subckt BUFT_X4_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE net_000 VSS N_ISO W=0.46e-06 L=0.18e-06
M1 VSS net_000 net_002 VSS N_ISO W=0.46e-06 L=0.18e-06
M2 net_002 OE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS net_002 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M6 VDD OE net_000 VDD P_ISO W=0.45e-06 L=0.18e-06
M7 VDD OE net_001 VDD P_ISO W=0.45e-06 L=0.18e-06
M8 net_001 net_000 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_001 A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD net_001 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M11 VDD net_001 Q VDD P_ISO W=1.05e-06 L=0.18e-06
.ends

.subckt BUFT_X6_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.71e-06 L=0.18e-06
M2 net_001 OE net_002 VSS N_ISO W=0.71e-06 L=0.18e-06
M3 VSS A net_001 VSS N_ISO W=0.71e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M7 VDD OE net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD OE net_002 VDD P_ISO W=0.78e-06 L=0.18e-06
M9 net_002 net_000 net_001 VDD P_ISO W=0.78e-06 L=0.18e-06
M10 VDD A net_002 VDD P_ISO W=0.755e-06 L=0.18e-06
M11 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M13 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
.ends

.subckt BUFT_X8_18_SVT_WB A OE Q VDD VSS
*.PININFO A:I OE:I Q:O VDD:B VSS:B
M0 VSS OE net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.71e-06 L=0.18e-06
M2 net_001 OE net_002 VSS N_ISO W=0.71e-06 L=0.18e-06
M3 VSS A net_001 VSS N_ISO W=0.71e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M7 VSS net_001 Q VSS N_ISO W=0.95e-06 L=0.18e-06
M8 VDD OE net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD OE net_002 VDD P_ISO W=0.78e-06 L=0.18e-06
M10 net_002 net_000 net_001 VDD P_ISO W=0.78e-06 L=0.18e-06
M11 VDD A net_002 VDD P_ISO W=0.755e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M13 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M15 VDD net_002 Q VDD P_ISO W=1.05e-06 L=0.18e-06
.ends

.subckt BUF_X10_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X12_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X14_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=0.815e-06 L=0.18e-06
M1 Q_neg A VSS VSS N_ISO W=0.815e-06 L=0.18e-06
M2 VSS A Q_neg VSS N_ISO W=0.815e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD A Q_neg VDD P_ISO W=0.895e-06 L=0.18e-06
M11 Q_neg A VDD VDD P_ISO W=0.895e-06 L=0.18e-06
M12 VDD A Q_neg VDD P_ISO W=0.895e-06 L=0.18e-06
M13 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X16_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X18_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X2_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VDD A Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M3 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X20_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X24_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X3_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=0.785e-06 L=0.18e-06
M1 Q Q_neg VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M2 VSS Q_neg Q VSS N_ISO W=0.785e-06 L=0.18e-06
M3 VDD A Q_neg VDD P_ISO W=0.86e-06 L=0.18e-06
M4 Q Q_neg VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M5 VDD Q_neg Q VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt BUF_X32_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.935e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=0.935e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=0.935e-06 L=0.18e-06
M3 VSS A net_000 VSS N_ISO W=0.935e-06 L=0.18e-06
M4 VSS A net_000 VSS N_ISO W=0.935e-06 L=0.18e-06
M5 VSS A net_000 VSS N_ISO W=0.935e-06 L=0.18e-06
M6 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VDD A net_000 VDD P_ISO W=1.02e-06 L=0.18e-06
M23 VDD A net_000 VDD P_ISO W=1.02e-06 L=0.18e-06
M24 VDD A net_000 VDD P_ISO W=1.02e-06 L=0.18e-06
M25 VDD A net_000 VDD P_ISO W=1.02e-06 L=0.18e-06
M26 VDD A net_000 VDD P_ISO W=1.02e-06 L=0.18e-06
M27 VDD A net_000 VDD P_ISO W=1.02e-06 L=0.18e-06
M28 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M42 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M4 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X5_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=0.58e-06 L=0.18e-06
.ends

.subckt BUF_X6_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M1 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A net_000 VDD P_ISO W=0.81e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt BUF_X8_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q_neg VSS N_ISO W=0.715e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q_neg A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A Q_neg VDD P_ISO W=0.815e-06 L=0.18e-06
M8 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKAND2_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.455e-06 L=0.18e-06
M1 net_001 A net_000 VSS N_ISO W=0.455e-06 L=0.18e-06
M2 net_001 A net_002 VSS N_ISO W=0.455e-06 L=0.18e-06
M3 VSS B net_002 VSS N_ISO W=0.455e-06 L=0.18e-06
M4 Q net_001 VSS VSS N_ISO W=0.455e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=0.455e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=0.45e-06 L=0.18e-06
M7 VSS net_001 Q VSS N_ISO W=0.45e-06 L=0.18e-06
M8 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q net_001 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_001 Q VDD P_ISO W=1.535e-06 L=0.18e-06
M14 VDD net_001 Q VDD P_ISO W=1.535e-06 L=0.18e-06
M15 VDD net_001 Q VDD P_ISO W=1.535e-06 L=0.18e-06
M16 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKAND2_X16_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_008 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_005 A net_008 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_009 A net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_010 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_005 A net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_011 A net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B net_011 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q net_005 VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M9 VSS net_005 Q VSS N_ISO W=0.475e-06 L=0.18e-06
M10 Q net_005 VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M11 VSS net_005 Q VSS N_ISO W=0.475e-06 L=0.18e-06
M12 Q net_005 VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M13 net_005 B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_005 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_005 B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_005 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 Q net_005 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M23 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M24 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M25 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M26 VDD net_005 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKAND2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.32e-06
M3 VDD A net_000 VDD P_ISO W=1.07e-06 L=0.18e-06
M4 VDD B net_000 VDD P_ISO W=1.07e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKAND2_X3_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 net_001 A net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 VSS net_001 Q VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD net_001 Q VDD P_ISO W=0.86e-06 L=0.18e-06
M6 VDD net_001 Q VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt CLKAND2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 net_001 A net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 VSS net_001 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M3 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKAND2_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 net_000 A net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 VSS net_001 Q VSS N_ISO W=0.915e-06 L=0.18e-06
M3 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKAND2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.455e-06 L=0.18e-06
M1 net_001 A net_000 VSS N_ISO W=0.455e-06 L=0.18e-06
M2 net_001 A net_002 VSS N_ISO W=0.455e-06 L=0.18e-06
M3 VSS B net_002 VSS N_ISO W=0.455e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M6 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X12_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.61e-06 L=0.18e-06
M1 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M2 Q net_000 VSS VSS N_ISO W=0.46e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M5 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M8 VDD net_000 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X16_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_004 A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS A net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q net_004 VSS VSS N_ISO W=0.495e-06 L=0.18e-06
M4 VSS net_004 Q VSS N_ISO W=0.495e-06 L=0.18e-06
M5 Q net_004 VSS VSS N_ISO W=0.495e-06 L=0.18e-06
M6 VSS net_004 Q VSS N_ISO W=0.495e-06 L=0.18e-06
M7 Q net_004 VSS VSS N_ISO W=0.495e-06 L=0.18e-06
M8 VDD A net_004 VDD P_ISO W=0.805e-06 L=0.18e-06
M9 net_004 A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M10 VDD A net_004 VDD P_ISO W=1.66e-06 L=0.18e-06
M11 Q net_004 VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M12 VDD net_004 Q VDD P_ISO W=1.61e-06 L=0.18e-06
M13 Q net_004 VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M14 VDD net_004 Q VDD P_ISO W=1.61e-06 L=0.18e-06
M15 Q net_004 VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M16 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X2_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 net_001 A VSS VSS N_ISO W=0.42e-06 L=0.23e-06
M1 Q net_001 VSS VSS N_ISO W=0.42e-06 L=0.23e-06
M2 net_001 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M3 Q net_001 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X20_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_005 VSS N_ISO W=0.475e-06 L=0.18e-06
M1 net_005 A VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M2 VSS A net_005 VSS N_ISO W=0.435e-06 L=0.18e-06
M3 Q net_005 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M4 VSS net_005 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M5 Q net_005 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M6 VSS net_005 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M7 Q net_005 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M8 VSS net_005 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M9 Q net_005 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M10 net_005 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A net_005 VDD P_ISO W=1.53e-06 L=0.18e-06
M12 net_005 A VDD VDD P_ISO W=1.53e-06 L=0.18e-06
M13 VDD A net_005 VDD P_ISO W=1.53e-06 L=0.18e-06
M14 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M15 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M16 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M17 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M18 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M19 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M20 Q net_005 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X24_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.46e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=0.46e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=0.46e-06 L=0.18e-06
M3 VSS A net_000 VSS N_ISO W=0.46e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M6 Q net_000 VSS VSS N_ISO W=0.46e-06 L=0.18e-06
M7 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M8 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M9 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M10 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M11 VSS net_000 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M12 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A net_000 VDD P_ISO W=1.44e-06 L=0.18e-06
M14 VDD A net_000 VDD P_ISO W=1.1e-06 L=0.18e-06
M15 VDD A net_000 VDD P_ISO W=1.44e-06 L=0.18e-06
M16 VDD A net_000 VDD P_ISO W=1.44e-06 L=0.18e-06
M17 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M18 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M19 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M20 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M21 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M22 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M23 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M24 VDD net_000 Q VDD P_ISO W=1.58e-06 L=0.18e-06
M25 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X3_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 net_001 A VSS VSS N_ISO W=0.42e-06 L=0.36e-06
M1 Q net_001 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_001 A VDD VDD P_ISO W=1.05e-06 L=0.18e-06
M3 Q net_001 VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M4 Q net_001 VDD VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt CLKBUF_X32_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_005 VSS N_ISO W=0.475e-06 L=0.18e-06
M1 net_005 A VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M2 VSS A net_005 VSS N_ISO W=0.475e-06 L=0.18e-06
M3 net_005 A VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M4 VSS A net_005 VSS N_ISO W=0.475e-06 L=0.18e-06
M5 Q net_005 VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M6 VSS net_005 Q VSS N_ISO W=0.445e-06 L=0.18e-06
M7 Q net_005 VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M8 VSS net_005 Q VSS N_ISO W=0.445e-06 L=0.18e-06
M9 Q net_005 VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M10 VSS net_005 Q VSS N_ISO W=0.445e-06 L=0.18e-06
M11 Q net_005 VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M12 VSS net_005 Q VSS N_ISO W=0.445e-06 L=0.18e-06
M13 Q net_005 VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M14 VSS net_005 Q VSS N_ISO W=0.445e-06 L=0.18e-06
M15 Q net_005 VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M16 net_005 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A net_005 VDD P_ISO W=1.61e-06 L=0.18e-06
M18 net_005 A VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M19 VDD A net_005 VDD P_ISO W=1.61e-06 L=0.18e-06
M20 net_005 A VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M21 VDD A net_005 VDD P_ISO W=1.61e-06 L=0.18e-06
M22 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M23 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M24 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M25 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M26 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M27 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M28 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M29 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M30 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M31 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M32 Q net_005 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 net_001 A VSS VSS N_ISO W=0.42e-06 L=0.36e-06
M1 Q net_001 VSS VSS N_ISO W=0.6e-06 L=0.18e-06
M2 net_001 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M3 Q net_001 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M4 Q net_001 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X40_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_004 VSS N_ISO W=0.435e-06 L=0.18e-06
M1 net_004 A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M2 VSS A net_004 VSS N_ISO W=0.435e-06 L=0.18e-06
M3 net_004 A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M4 VSS A net_004 VSS N_ISO W=0.435e-06 L=0.18e-06
M5 net_004 A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M6 VSS A net_004 VSS N_ISO W=0.435e-06 L=0.18e-06
M7 Q net_004 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M8 VSS net_004 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M9 Q net_004 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M10 VSS net_004 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M11 Q net_004 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M12 VSS net_004 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M13 Q net_004 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M14 VSS net_004 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M15 Q net_004 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M16 VSS net_004 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M17 Q net_004 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M18 VSS net_004 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M19 Q net_004 VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M20 VSS net_004 Q VSS N_ISO W=0.435e-06 L=0.18e-06
M21 VDD A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_004 A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M23 VDD A net_004 VDD P_ISO W=1.66e-06 L=0.18e-06
M24 net_004 A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M25 VDD A net_004 VDD P_ISO W=1.66e-06 L=0.18e-06
M26 net_004 A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M27 VDD A net_004 VDD P_ISO W=1.66e-06 L=0.18e-06
M28 Q net_004 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M29 VDD net_004 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M30 Q net_004 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M31 VDD net_004 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M32 Q net_004 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M33 VDD net_004 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M34 Q net_004 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M35 VDD net_004 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M36 Q net_004 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M37 VDD net_004 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M38 Q net_004 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M39 VDD net_004 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M40 Q net_004 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M41 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKBUF_X6_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q net_004 VSS VSS N_ISO W=0.46e-06 L=0.18e-06
M2 VSS net_004 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M3 VDD A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 Q net_004 VDD VDD P_ISO W=1.32e-06 L=0.18e-06
M5 VDD net_004 Q VDD P_ISO W=1.66e-06 L=0.18e-06
.ends

.subckt CLKBUF_X8_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_005 VSS N_ISO W=0.465e-06 L=0.18e-06
M1 Q net_005 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_005 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q net_005 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_005 A VDD VDD P_ISO W=0.81e-06 L=0.18e-06
M5 VDD A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q net_005 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M7 VDD net_005 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M8 Q net_005 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X1_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.42e-06 L=0.44e-06
M1 Q A VDD VDD P_ISO W=0.9e-06 L=0.18e-06
.ends

.subckt CLKINV_X12_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.45e-06 L=0.18e-06
M1 Q A VSS VSS N_ISO W=0.45e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.45e-06 L=0.18e-06
M3 Q A VSS VSS N_ISO W=0.45e-06 L=0.18e-06
M4 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q A VDD VDD P_ISO W=1.535e-06 L=0.18e-06
M6 Q A VDD VDD P_ISO W=1.535e-06 L=0.18e-06
M7 Q A VDD VDD P_ISO W=1.535e-06 L=0.18e-06
M8 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X16_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.475e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.475e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M5 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M7 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M9 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X2_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.42e-06 L=0.32e-06
M1 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X20_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M7 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.535e-06 L=0.18e-06
M9 Q A VDD VDD P_ISO W=1.535e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.535e-06 L=0.18e-06
M11 Q A VDD VDD P_ISO W=1.535e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.535e-06 L=0.18e-06
M13 Q A VDD VDD P_ISO W=1.535e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X24_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.46e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.46e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.46e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.46e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.46e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.46e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=0.46e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.46e-06 L=0.18e-06
M8 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.645e-06 L=0.18e-06
M10 Q A VDD VDD P_ISO W=1.645e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.645e-06 L=0.18e-06
M12 Q A VDD VDD P_ISO W=1.645e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.645e-06 L=0.18e-06
M14 Q A VDD VDD P_ISO W=1.645e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.645e-06 L=0.18e-06
M16 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X3_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.44e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt CLKINV_X32_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.445e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.445e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.445e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.445e-06 L=0.18e-06
M8 Q A VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.445e-06 L=0.18e-06
M10 Q A VSS VSS N_ISO W=0.445e-06 L=0.18e-06
M11 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.61e-06 L=0.18e-06
M13 Q A VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.61e-06 L=0.18e-06
M15 Q A VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.61e-06 L=0.18e-06
M17 Q A VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=1.61e-06 L=0.18e-06
M19 Q A VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M20 VDD A Q VDD P_ISO W=1.61e-06 L=0.18e-06
M21 Q A VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M22 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.61e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X40_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M8 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M10 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M12 Q A VSS VSS N_ISO W=0.435e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=0.435e-06 L=0.18e-06
M14 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M16 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M18 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M19 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M20 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M22 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M23 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M24 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M26 Q A VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M27 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X6_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.915e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M3 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKINV_X8_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.61e-06 L=0.18e-06
M1 Q A VSS VSS N_ISO W=0.61e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M3 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M4 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKMUX2_X12_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_004 net_005 VSS N_ISO W=0.915e-06 L=0.18e-06
M7 VSS net_005 Q VSS N_ISO W=0.45e-06 L=0.18e-06
M8 VSS net_005 Q VSS N_ISO W=0.45e-06 L=0.18e-06
M9 VSS net_005 Q VSS N_ISO W=0.45e-06 L=0.18e-06
M10 VSS net_005 Q VSS N_ISO W=0.45e-06 L=0.18e-06
M11 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD B net_006 VDD P_ISO W=0.865e-06 L=0.18e-06
M13 net_002 net_000 net_006 VDD P_ISO W=0.865e-06 L=0.18e-06
M14 net_002 S0 net_007 VDD P_ISO W=0.865e-06 L=0.18e-06
M15 VDD A net_007 VDD P_ISO W=0.865e-06 L=0.18e-06
M16 VDD net_002 net_004 VDD P_ISO W=0.865e-06 L=0.18e-06
M17 VDD net_002 net_004 VDD P_ISO W=0.865e-06 L=0.18e-06
M18 VDD net_004 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_004 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_004 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_005 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_005 Q VDD P_ISO W=1.535e-06 L=0.18e-06
M23 VDD net_005 Q VDD P_ISO W=1.535e-06 L=0.18e-06
M24 VDD net_005 Q VDD P_ISO W=1.535e-06 L=0.18e-06
M25 VDD net_005 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKMUX2_X16_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_012 B VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_007 S0 net_012 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_013 net_004 net_007 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_013 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_009 net_007 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_007 net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_010 net_009 VSS VSS N_ISO W=0.61e-06 L=0.18e-06
M8 VSS net_009 net_010 VSS N_ISO W=0.61e-06 L=0.18e-06
M9 Q net_010 VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M10 VSS net_010 Q VSS N_ISO W=0.475e-06 L=0.18e-06
M11 Q net_010 VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M12 VSS net_010 Q VSS N_ISO W=0.475e-06 L=0.18e-06
M13 Q net_010 VSS VSS N_ISO W=0.475e-06 L=0.18e-06
M14 VDD S0 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M15 net_014 B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M16 net_007 net_004 net_014 VDD P_ISO W=0.575e-06 L=0.18e-06
M17 net_015 S0 net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M18 VDD A net_015 VDD P_ISO W=0.575e-06 L=0.18e-06
M19 net_009 net_007 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_007 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_010 net_009 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_009 net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 net_010 net_009 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_009 net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M25 Q net_010 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_010 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M27 Q net_010 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=1.66e-06 L=0.18e-06
M29 Q net_010 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M30 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKMUX2_X2_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.45e-06 L=0.18e-06
M6 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_002 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_002 S0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKMUX2_X3_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B net_004 VDD P_ISO W=0.865e-06 L=0.18e-06
M8 net_002 net_000 net_004 VDD P_ISO W=0.865e-06 L=0.18e-06
M9 net_002 S0 net_005 VDD P_ISO W=0.865e-06 L=0.18e-06
M10 VDD A net_005 VDD P_ISO W=0.865e-06 L=0.18e-06
M11 VDD net_002 Q VDD P_ISO W=0.865e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=0.865e-06 L=0.18e-06
.ends

.subckt CLKMUX2_X4_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_002 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_002 S0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKMUX2_X6_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.915e-06 L=0.18e-06
M6 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_002 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_002 S0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKMUX2_X8_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M7 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_002 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_005 S0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_005 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKNAND2_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.535e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=0.535e-06 L=0.18e-06
M2 net_001 A Q VSS N_ISO W=0.535e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=0.535e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=0.535e-06 L=0.18e-06
M5 Q A net_002 VSS N_ISO W=0.535e-06 L=0.18e-06
M6 Q A net_003 VSS N_ISO W=0.535e-06 L=0.18e-06
M7 VSS B net_003 VSS N_ISO W=0.535e-06 L=0.18e-06
M8 VSS B net_004 VSS N_ISO W=0.535e-06 L=0.18e-06
M9 Q A net_004 VSS N_ISO W=0.535e-06 L=0.18e-06
M10 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.44e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.44e-06 L=0.18e-06
M13 VDD B Q VDD P_ISO W=1.44e-06 L=0.18e-06
M14 VDD B Q VDD P_ISO W=1.44e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.44e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.44e-06 L=0.18e-06
M17 VDD B Q VDD P_ISO W=1.44e-06 L=0.18e-06
M18 VDD B Q VDD P_ISO W=1.44e-06 L=0.18e-06
M19 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKNAND2_X16_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.51e-06 L=0.18e-06
M1 Q B net_000 VSS N_ISO W=0.51e-06 L=0.18e-06
M2 Q B net_001 VSS N_ISO W=0.51e-06 L=0.18e-06
M3 VSS A net_001 VSS N_ISO W=0.51e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=0.51e-06 L=0.18e-06
M5 Q B net_002 VSS N_ISO W=0.51e-06 L=0.18e-06
M6 net_003 B Q VSS N_ISO W=0.51e-06 L=0.18e-06
M7 VSS A net_003 VSS N_ISO W=0.51e-06 L=0.18e-06
M8 VSS A net_004 VSS N_ISO W=0.51e-06 L=0.18e-06
M9 Q B net_004 VSS N_ISO W=0.51e-06 L=0.18e-06
M10 Q B net_005 VSS N_ISO W=0.51e-06 L=0.18e-06
M11 VSS A net_005 VSS N_ISO W=0.51e-06 L=0.18e-06
M12 VSS A net_006 VSS N_ISO W=0.51e-06 L=0.18e-06
M13 Q B net_006 VSS N_ISO W=0.51e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.34e-06 L=0.18e-06
M16 VDD B Q VDD P_ISO W=1.34e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.34e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=1.34e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=1.34e-06 L=0.18e-06
M20 VDD B Q VDD P_ISO W=1.34e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.34e-06 L=0.18e-06
M22 VDD A Q VDD P_ISO W=1.34e-06 L=0.18e-06
M23 VDD B Q VDD P_ISO W=1.34e-06 L=0.18e-06
M24 VDD B Q VDD P_ISO W=1.34e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.34e-06 L=0.18e-06
M26 VDD A Q VDD P_ISO W=1.34e-06 L=0.18e-06
M27 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKNAND2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKNAND2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.455e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=0.455e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=0.455e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=0.455e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKNAND2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M5 Q A net_002 VSS N_ISO W=0.45e-06 L=0.18e-06
M6 Q A net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M7 VSS B net_003 VSS N_ISO W=0.45e-06 L=0.18e-06
M8 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKXOR2_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_003 A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_003 B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_003 net_004 VSS N_ISO W=0.61e-06 L=0.18e-06
M6 VSS net_004 net_005 VSS N_ISO W=0.61e-06 L=0.18e-06
M7 VSS net_005 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M8 VSS net_005 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M9 VSS net_005 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M10 VSS net_005 Q VSS N_ISO W=0.46e-06 L=0.18e-06
M11 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_003 A net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_003 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_003 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_004 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_004 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_005 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M21 VDD net_005 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M22 VDD net_005 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M23 VDD net_005 Q VDD P_ISO W=1.44e-06 L=0.18e-06
M24 VDD net_005 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKXOR2_X16_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_012 A net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_012 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_007 net_004 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_008 A net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_007 B net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_009 net_008 VSS VSS N_ISO W=0.61e-06 L=0.18e-06
M6 VSS net_008 net_009 VSS N_ISO W=0.61e-06 L=0.18e-06
M7 VSS net_009 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_010 net_009 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M9 VSS net_009 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 Q net_010 VSS VSS N_ISO W=0.495e-06 L=0.18e-06
M11 VSS net_010 Q VSS N_ISO W=0.495e-06 L=0.18e-06
M12 Q net_010 VSS VSS N_ISO W=0.495e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.495e-06 L=0.18e-06
M14 Q net_010 VSS VSS N_ISO W=0.495e-06 L=0.18e-06
M15 net_004 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_008 net_004 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_013 A net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B net_013 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 net_009 net_008 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_008 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_009 net_008 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_008 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_009 net_010 VDD P_ISO W=0.805e-06 L=0.18e-06
M25 net_010 net_009 VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M26 VDD net_009 net_010 VDD P_ISO W=1.66e-06 L=0.18e-06
M27 Q net_010 VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=1.61e-06 L=0.18e-06
M29 Q net_010 VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M30 VDD net_010 Q VDD P_ISO W=1.61e-06 L=0.18e-06
M31 Q net_010 VDD VDD P_ISO W=1.61e-06 L=0.18e-06
M32 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKXOR2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_002 A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKXOR2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_003 A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_003 B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_003 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M6 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_003 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt CLKXOR2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_003 A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_003 B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_003 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=0.61e-06 L=0.18e-06
M7 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_003 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFQN_X1_18_SVT_WB D CK QN VDD VSS
*.PININFO D:I CK:I QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.425e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS net_006 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M12 VDD CK net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M13 VDD net_000 net_001 VDD P_ISO W=0.725e-06 L=0.18e-06
M14 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M15 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M16 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M17 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 VDD net_003 net_005 VDD P_ISO W=0.435e-06 L=0.18e-06
M19 net_006 net_000 net_005 VDD P_ISO W=0.56e-06 L=0.18e-06
M20 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_006 net_008 VDD P_ISO W=0.415e-06 L=0.18e-06
M23 VDD net_006 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFFQN_X2_18_SVT_WB D CK QN VDD VSS
*.PININFO D:I CK:I QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.52e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS net_006 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M12 VDD CK net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M13 VDD net_000 net_001 VDD P_ISO W=0.725e-06 L=0.18e-06
M14 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M15 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M16 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M17 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 VDD net_003 net_005 VDD P_ISO W=0.685e-06 L=0.18e-06
M19 net_006 net_000 net_005 VDD P_ISO W=0.71e-06 L=0.18e-06
M20 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_006 net_008 VDD P_ISO W=0.415e-06 L=0.18e-06
M23 VDD net_006 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFQN_X4_18_SVT_WB D CK QN VDD VSS
*.PININFO D:I CK:I QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS net_006 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M12 VSS net_006 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M13 VDD CK net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M14 VDD net_000 net_001 VDD P_ISO W=0.725e-06 L=0.18e-06
M15 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M16 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M17 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M19 VDD net_003 net_005 VDD P_ISO W=0.685e-06 L=0.18e-06
M20 net_006 net_000 net_005 VDD P_ISO W=0.755e-06 L=0.18e-06
M21 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M23 VDD net_006 net_008 VDD P_ISO W=0.415e-06 L=0.18e-06
M24 VDD net_006 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_006 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFQ_X1_18_SVT_WB D CK Q VDD VSS
*.PININFO D:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M12 VDD CK net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M13 VDD net_000 net_001 VDD P_ISO W=0.725e-06 L=0.18e-06
M14 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M15 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M16 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M17 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 net_005 net_003 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M19 net_006 net_000 net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_006 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_008 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFFQ_X2_18_SVT_WB D CK Q VDD VSS
*.PININFO D:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.535e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M12 VDD CK net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M13 VDD net_000 net_001 VDD P_ISO W=0.725e-06 L=0.18e-06
M14 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M15 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M16 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M17 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 net_005 net_003 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M19 net_006 net_000 net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_006 net_008 VDD P_ISO W=0.59e-06 L=0.18e-06
M23 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFQ_X4_18_SVT_WB D CK Q VDD VSS
*.PININFO D:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_005 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.535e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M12 VSS net_008 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M13 VDD CK net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M14 VDD net_000 net_001 VDD P_ISO W=0.725e-06 L=0.18e-06
M15 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M16 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M17 net_003 net_000 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 VDD net_005 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 net_005 net_003 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M20 net_006 net_000 net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 net_006 net_001 net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_008 net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_006 net_008 VDD P_ISO W=0.59e-06 L=0.18e-06
M24 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFQ_X8_18_SVT_WB D CK Q VDD VSS
*.PININFO D:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.535e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M12 VSS net_008 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M13 VSS net_008 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M14 VSS net_008 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.725e-06 L=0.18e-06
M17 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M18 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M19 net_003 net_000 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD net_005 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 net_005 net_003 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M22 net_006 net_000 net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 net_006 net_001 net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_008 net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_006 net_008 VDD P_ISO W=0.59e-06 L=0.18e-06
M26 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFRQ_X1_18_SVT_WB D RN CK Q VDD VSS
*.PININFO D:I RN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.55e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.475e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 net_005 RN net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_007 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_010 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS RN net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 net_007 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M14 VDD CK net_000 VDD P_ISO W=0.48e-06 L=0.18e-06
M15 VDD net_000 net_001 VDD P_ISO W=0.62e-06 L=0.18e-06
M16 VDD net_001 net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M17 net_003 D net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M18 net_003 net_000 net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD RN net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD net_006 net_012 VDD P_ISO W=0.425e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=0.53e-06 L=0.18e-06
M22 net_007 net_000 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 net_007 net_001 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M24 VDD net_010 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD RN net_010 VDD P_ISO W=0.415e-06 L=0.18e-06
M26 VDD net_007 net_010 VDD P_ISO W=0.545e-06 L=0.18e-06
M27 VDD net_010 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFFRQ_X2_18_SVT_WB D RN CK Q VDD VSS
*.PININFO D:I RN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.53e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 net_005 RN net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.51e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_007 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_010 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS RN net_009 VSS N_ISO W=0.495e-06 L=0.18e-06
M12 net_010 net_007 net_009 VSS N_ISO W=0.495e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M14 VDD CK net_000 VDD P_ISO W=0.505e-06 L=0.18e-06
M15 VDD net_000 net_001 VDD P_ISO W=0.745e-06 L=0.18e-06
M16 VDD net_001 net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M17 net_003 D net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M18 net_003 net_000 net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD RN net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD net_006 net_012 VDD P_ISO W=0.425e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=0.685e-06 L=0.18e-06
M22 net_007 net_000 net_006 VDD P_ISO W=0.545e-06 L=0.18e-06
M23 net_007 net_001 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M24 VDD net_010 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD RN net_010 VDD P_ISO W=0.415e-06 L=0.18e-06
M26 VDD net_007 net_010 VDD P_ISO W=0.715e-06 L=0.18e-06
M27 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFRQ_X4_18_SVT_WB D RN CK Q VDD VSS
*.PININFO D:I RN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.56e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.465e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 net_005 RN net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 net_006 net_003 VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_007 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_010 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS RN net_009 VSS N_ISO W=0.525e-06 L=0.18e-06
M12 net_010 net_007 net_009 VSS N_ISO W=0.525e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.47e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.62e-06 L=0.18e-06
M17 VDD net_001 net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M18 net_003 D net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M19 net_012 net_000 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD RN net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD net_006 net_012 VDD P_ISO W=0.425e-06 L=0.18e-06
M22 VDD net_003 net_006 VDD P_ISO W=0.65e-06 L=0.18e-06
M23 net_007 net_000 net_006 VDD P_ISO W=0.495e-06 L=0.18e-06
M24 net_007 net_001 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_010 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD RN net_010 VDD P_ISO W=0.415e-06 L=0.18e-06
M27 VDD net_007 net_010 VDD P_ISO W=0.715e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFRQ_X8_18_SVT_WB D RN CK Q VDD VSS
*.PININFO D:I RN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.56e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.465e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 net_005 RN net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.695e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.57e-06 L=0.18e-06
M9 net_007 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_010 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS RN net_009 VSS N_ISO W=0.925e-06 L=0.18e-06
M12 net_010 net_007 net_009 VSS N_ISO W=0.925e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M15 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M16 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.47e-06 L=0.18e-06
M18 VDD net_000 net_001 VDD P_ISO W=0.62e-06 L=0.18e-06
M19 VDD net_001 net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M20 net_003 D net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M21 net_003 net_000 net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD RN net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_006 net_012 VDD P_ISO W=0.425e-06 L=0.18e-06
M24 VDD net_003 net_006 VDD P_ISO W=0.71e-06 L=0.18e-06
M25 net_007 net_000 net_006 VDD P_ISO W=0.675e-06 L=0.18e-06
M26 net_007 net_001 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_010 net_013 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD RN net_010 VDD P_ISO W=0.415e-06 L=0.18e-06
M29 VDD net_007 net_010 VDD P_ISO W=1.145e-06 L=0.18e-06
M30 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFR_X1_18_SVT_WB D RN CK Q QN VDD VSS
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.535e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.465e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 net_005 RN net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_010 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS RN net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 net_007 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M14 VSS net_008 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.465e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.61e-06 L=0.18e-06
M17 VDD net_001 net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M18 net_003 D net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M19 net_003 net_000 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 VDD RN net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD net_006 net_012 VDD P_ISO W=0.425e-06 L=0.18e-06
M22 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 net_007 net_000 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_008 net_001 net_007 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_010 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD RN net_010 VDD P_ISO W=0.415e-06 L=0.18e-06
M27 VDD net_007 net_010 VDD P_ISO W=0.625e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M29 VDD net_008 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFFR_X2_18_SVT_WB D RN CK Q QN VDD VSS
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.435e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 net_005 RN net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_010 net_008 VSS N_ISO W=0.56e-06 L=0.18e-06
M11 VSS RN net_009 VSS N_ISO W=0.56e-06 L=0.18e-06
M12 net_010 net_007 net_009 VSS N_ISO W=0.56e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M14 VSS net_008 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.5e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.645e-06 L=0.18e-06
M17 VDD net_001 net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M18 net_003 D net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M19 net_012 net_000 net_003 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 VDD RN net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD net_006 net_012 VDD P_ISO W=0.425e-06 L=0.18e-06
M22 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 net_007 net_000 net_006 VDD P_ISO W=0.595e-06 L=0.18e-06
M24 net_008 net_001 net_007 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_010 net_008 VDD P_ISO W=0.67e-06 L=0.18e-06
M26 VDD RN net_010 VDD P_ISO W=0.415e-06 L=0.18e-06
M27 VDD net_007 net_010 VDD P_ISO W=0.715e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFR_X4_18_SVT_WB D RN CK Q QN VDD VSS
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 net_005 RN net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.545e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.49e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_010 net_008 VSS N_ISO W=0.7e-06 L=0.18e-06
M11 VSS RN net_009 VSS N_ISO W=0.7e-06 L=0.18e-06
M12 net_010 net_007 net_009 VSS N_ISO W=0.7e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M15 VSS net_008 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M16 VSS net_008 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.495e-06 L=0.18e-06
M18 VDD net_000 net_001 VDD P_ISO W=0.76e-06 L=0.18e-06
M19 VDD net_001 net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M20 net_003 D net_011 VDD P_ISO W=0.685e-06 L=0.18e-06
M21 net_003 net_000 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD RN net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 net_012 net_006 VDD VDD P_ISO W=0.425e-06 L=0.18e-06
M24 VDD net_003 net_006 VDD P_ISO W=0.57e-06 L=0.18e-06
M25 net_007 net_000 net_006 VDD P_ISO W=0.545e-06 L=0.18e-06
M26 net_008 net_001 net_007 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 net_008 net_010 VDD VDD P_ISO W=0.655e-06 L=0.18e-06
M28 VDD RN net_010 VDD P_ISO W=0.415e-06 L=0.18e-06
M29 VDD net_007 net_010 VDD P_ISO W=0.715e-06 L=0.18e-06
M30 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFS_PX8_18_SVT_WB D SN CK Q QN VDD VSS
*.PININFO D:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.59e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.82e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.82e-06 L=0.18e-06
M8 net_006 net_001 net_007 VSS N_ISO W=0.545e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.84e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.67e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_007 net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M24 VDD net_001 net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M25 net_003 D net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M26 net_003 net_000 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_006 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_003 net_006 VDD P_ISO W=1.015e-06 L=0.18e-06
M29 VDD SN net_006 VDD P_ISO W=0.45e-06 L=0.18e-06
M30 net_007 net_000 net_006 VDD P_ISO W=0.74e-06 L=0.18e-06
M31 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M32 VDD SN net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M33 VDD net_010 net_008 VDD P_ISO W=0.815e-06 L=0.18e-06
M34 VDD net_007 net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD net_007 net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M42 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFSQ_X1_18_SVT_WB D SN CK Q VDD VSS
*.PININFO D:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.475e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.505e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=0.44e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M14 VDD CK net_000 VDD P_ISO W=0.5e-06 L=0.18e-06
M15 VDD net_000 net_001 VDD P_ISO W=0.675e-06 L=0.18e-06
M16 VDD net_001 net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M17 net_003 D net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M18 net_003 net_000 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M19 VDD net_006 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M20 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SN net_006 VDD P_ISO W=0.655e-06 L=0.18e-06
M22 net_007 net_000 net_006 VDD P_ISO W=0.73e-06 L=0.18e-06
M23 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD SN net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 VDD net_010 net_008 VDD P_ISO W=0.45e-06 L=0.18e-06
M26 VDD net_007 net_010 VDD P_ISO W=0.455e-06 L=0.18e-06
M27 VDD net_010 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFFSQ_X2_18_SVT_WB D SN CK Q VDD VSS
*.PININFO D:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.475e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.505e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=0.62e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD CK net_000 VDD P_ISO W=0.5e-06 L=0.18e-06
M15 VDD net_000 net_001 VDD P_ISO W=0.675e-06 L=0.18e-06
M16 VDD net_001 net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M17 net_003 D net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M18 net_003 net_000 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M19 VDD net_006 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M20 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SN net_006 VDD P_ISO W=0.655e-06 L=0.18e-06
M22 net_007 net_000 net_006 VDD P_ISO W=0.73e-06 L=0.18e-06
M23 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD SN net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 VDD net_010 net_008 VDD P_ISO W=0.45e-06 L=0.18e-06
M26 VDD net_007 net_010 VDD P_ISO W=0.68e-06 L=0.18e-06
M27 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFSQ_X4_18_SVT_WB D SN CK Q VDD VSS
*.PININFO D:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.475e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.505e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=0.62e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.5e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.675e-06 L=0.18e-06
M17 VDD net_001 net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M18 net_003 D net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M19 net_003 net_000 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M20 VDD net_006 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD SN net_006 VDD P_ISO W=0.655e-06 L=0.18e-06
M23 net_007 net_000 net_006 VDD P_ISO W=0.73e-06 L=0.18e-06
M24 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD SN net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M26 VDD net_010 net_008 VDD P_ISO W=0.45e-06 L=0.18e-06
M27 VDD net_007 net_010 VDD P_ISO W=0.68e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFSQ_X8_18_SVT_WB D SN CK Q VDD VSS
*.PININFO D:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.475e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.505e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.505e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.675e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=0.62e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.5e-06 L=0.18e-06
M18 VDD net_000 net_001 VDD P_ISO W=0.675e-06 L=0.18e-06
M19 VDD net_001 net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M20 net_003 D net_011 VDD P_ISO W=0.6e-06 L=0.18e-06
M21 net_003 net_000 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M22 VDD net_006 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M23 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD SN net_006 VDD P_ISO W=0.655e-06 L=0.18e-06
M25 net_007 net_000 net_006 VDD P_ISO W=0.73e-06 L=0.18e-06
M26 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD SN net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M28 VDD net_010 net_008 VDD P_ISO W=0.45e-06 L=0.18e-06
M29 VDD net_007 net_010 VDD P_ISO W=0.68e-06 L=0.18e-06
M30 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFSR_X1_18_SVT_WB D RN SN CK Q QN VDD VSS
*.PININFO D:I RN:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 D VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_004 net_001 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_004 net_007 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 net_008 net_001 net_007 VSS N_ISO W=0.49e-06 L=0.18e-06
M10 net_009 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 net_009 SN net_010 VSS N_ISO W=0.62e-06 L=0.18e-06
M12 VSS net_012 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 VSS RN net_011 VSS N_ISO W=0.825e-06 L=0.18e-06
M14 net_011 net_008 net_012 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 VSS net_012 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M16 VSS net_009 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.45e-06 L=0.18e-06
M18 VDD net_000 net_001 VDD P_ISO W=0.76e-06 L=0.18e-06
M19 VDD D net_002 VDD P_ISO W=0.585e-06 L=0.18e-06
M20 net_003 net_001 net_002 VDD P_ISO W=0.585e-06 L=0.18e-06
M21 net_003 net_000 net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M22 VDD net_007 net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M23 VDD RN net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M24 VDD net_003 net_007 VDD P_ISO W=0.45e-06 L=0.18e-06
M25 VDD SN net_007 VDD P_ISO W=0.45e-06 L=0.18e-06
M26 net_008 net_000 net_007 VDD P_ISO W=0.585e-06 L=0.18e-06
M27 net_008 net_001 net_009 VDD P_ISO W=0.45e-06 L=0.18e-06
M28 VDD SN net_009 VDD P_ISO W=0.625e-06 L=0.18e-06
M29 VDD net_012 net_009 VDD P_ISO W=0.815e-06 L=0.18e-06
M30 VDD RN net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M31 VDD net_008 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M32 VDD net_012 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M33 VDD net_009 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFFSR_X2_18_SVT_WB D RN SN CK Q QN VDD VSS
*.PININFO D:I RN:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 D VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_004 net_001 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_004 net_007 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 net_008 net_001 net_007 VSS N_ISO W=0.49e-06 L=0.18e-06
M10 net_009 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 net_009 SN net_010 VSS N_ISO W=0.62e-06 L=0.18e-06
M12 VSS net_012 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 VSS RN net_011 VSS N_ISO W=0.825e-06 L=0.18e-06
M14 net_011 net_008 net_012 VSS N_ISO W=0.92e-06 L=0.18e-06
M15 VSS net_012 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_009 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.45e-06 L=0.18e-06
M18 VDD net_000 net_001 VDD P_ISO W=0.76e-06 L=0.18e-06
M19 VDD D net_002 VDD P_ISO W=0.585e-06 L=0.18e-06
M20 net_003 net_001 net_002 VDD P_ISO W=0.585e-06 L=0.18e-06
M21 net_003 net_000 net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M22 VDD net_007 net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M23 VDD RN net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M24 VDD net_003 net_007 VDD P_ISO W=0.45e-06 L=0.18e-06
M25 VDD SN net_007 VDD P_ISO W=0.45e-06 L=0.18e-06
M26 net_008 net_000 net_007 VDD P_ISO W=0.585e-06 L=0.18e-06
M27 net_008 net_001 net_009 VDD P_ISO W=0.45e-06 L=0.18e-06
M28 VDD SN net_009 VDD P_ISO W=0.625e-06 L=0.18e-06
M29 VDD net_012 net_009 VDD P_ISO W=0.815e-06 L=0.18e-06
M30 VDD RN net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M31 VDD net_008 net_012 VDD P_ISO W=0.96e-06 L=0.18e-06
M32 VDD net_012 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_009 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFSR_X4_18_SVT_WB D RN SN CK Q QN VDD VSS
*.PININFO D:I RN:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.62e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 D VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_004 net_001 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_004 net_007 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 net_008 net_001 net_007 VSS N_ISO W=0.49e-06 L=0.18e-06
M10 net_009 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 net_009 SN net_010 VSS N_ISO W=0.62e-06 L=0.18e-06
M12 VSS net_012 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 VSS RN net_011 VSS N_ISO W=0.825e-06 L=0.18e-06
M14 net_011 net_008 net_012 VSS N_ISO W=0.92e-06 L=0.18e-06
M15 VSS net_012 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_012 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_009 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_009 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.45e-06 L=0.18e-06
M20 VDD net_000 net_001 VDD P_ISO W=0.76e-06 L=0.18e-06
M21 VDD D net_002 VDD P_ISO W=0.585e-06 L=0.18e-06
M22 net_003 net_001 net_002 VDD P_ISO W=0.585e-06 L=0.18e-06
M23 net_003 net_000 net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M24 VDD net_007 net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M25 VDD RN net_013 VDD P_ISO W=0.45e-06 L=0.18e-06
M26 VDD net_003 net_007 VDD P_ISO W=0.45e-06 L=0.18e-06
M27 VDD SN net_007 VDD P_ISO W=0.45e-06 L=0.18e-06
M28 net_008 net_000 net_007 VDD P_ISO W=0.585e-06 L=0.18e-06
M29 net_008 net_001 net_009 VDD P_ISO W=0.45e-06 L=0.18e-06
M30 VDD SN net_009 VDD P_ISO W=0.625e-06 L=0.18e-06
M31 VDD net_012 net_009 VDD P_ISO W=0.815e-06 L=0.18e-06
M32 VDD RN net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M33 VDD net_008 net_012 VDD P_ISO W=0.96e-06 L=0.18e-06
M34 VDD net_012 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD net_012 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_009 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_009 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFS_X1_18_SVT_WB D SN CK Q QN VDD VSS
*.PININFO D:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.59e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.545e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.79e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.79e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M14 VSS net_008 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M17 VDD net_001 net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M18 net_003 D net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M19 net_003 net_000 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 VDD net_006 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD SN net_006 VDD P_ISO W=0.64e-06 L=0.18e-06
M23 net_007 net_000 net_006 VDD P_ISO W=0.695e-06 L=0.18e-06
M24 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD SN net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_010 net_008 VDD P_ISO W=0.84e-06 L=0.18e-06
M27 VDD net_007 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M29 VDD net_008 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFFS_X2_18_SVT_WB D SN CK Q QN VDD VSS
*.PININFO D:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.59e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.545e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.79e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.79e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=1.005e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M17 VDD net_001 net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M18 net_003 D net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M19 net_003 net_000 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 VDD net_006 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD SN net_006 VDD P_ISO W=0.64e-06 L=0.18e-06
M23 net_007 net_000 net_006 VDD P_ISO W=0.695e-06 L=0.18e-06
M24 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD SN net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_010 net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_007 net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFS_X4_18_SVT_WB D SN CK Q QN VDD VSS
*.PININFO D:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.59e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.545e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.79e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.79e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=1.005e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M19 VDD net_001 net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M20 net_003 D net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M21 net_003 net_000 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_006 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M23 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD SN net_006 VDD P_ISO W=0.64e-06 L=0.18e-06
M25 net_007 net_000 net_006 VDD P_ISO W=0.695e-06 L=0.18e-06
M26 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD SN net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M28 VDD net_010 net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_007 net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFS_X8_18_SVT_WB D SN CK Q QN VDD VSS
*.PININFO D:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.59e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.585e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_006 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M7 net_006 SN net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.545e-06 L=0.18e-06
M9 net_008 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 net_008 SN net_009 VSS N_ISO W=0.84e-06 L=0.18e-06
M11 VSS net_010 net_009 VSS N_ISO W=0.625e-06 L=0.18e-06
M12 VSS net_007 net_010 VSS N_ISO W=1.005e-06 L=0.18e-06
M13 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_010 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_008 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M23 VDD net_001 net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M24 net_003 D net_011 VDD P_ISO W=0.57e-06 L=0.18e-06
M25 net_003 net_000 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_006 net_012 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M28 VDD SN net_006 VDD P_ISO W=0.64e-06 L=0.18e-06
M29 net_007 net_000 net_006 VDD P_ISO W=0.695e-06 L=0.18e-06
M30 net_007 net_001 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M31 VDD SN net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M32 VDD net_010 net_008 VDD P_ISO W=0.815e-06 L=0.18e-06
M33 VDD net_007 net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_010 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_008 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFTR_X1_18_SVT_WB D RN CK Q QN VDD VSS
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.66e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 VSS RN net_002 VSS N_ISO W=0.54e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.54e-06 L=0.18e-06
M4 net_004 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M5 net_004 net_001 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_004 net_006 VSS N_ISO W=0.565e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_007 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_007 net_009 VSS N_ISO W=0.525e-06 L=0.18e-06
M13 VSS net_009 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M15 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M16 VDD RN net_003 VDD P_ISO W=0.475e-06 L=0.18e-06
M17 VDD D net_003 VDD P_ISO W=0.72e-06 L=0.18e-06
M18 net_004 net_001 net_003 VDD P_ISO W=0.41e-06 L=0.18e-06
M19 net_004 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 VDD net_006 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_004 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 net_007 net_000 net_006 VDD P_ISO W=0.565e-06 L=0.18e-06
M23 net_007 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M24 VDD net_009 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_007 net_009 VDD P_ISO W=0.575e-06 L=0.18e-06
M27 VDD net_009 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFTR_X2_18_SVT_WB D RN CK Q QN VDD VSS
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.66e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 VSS RN net_002 VSS N_ISO W=0.54e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.54e-06 L=0.18e-06
M4 net_004 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M5 net_004 net_001 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_004 net_006 VSS N_ISO W=0.59e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_007 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_007 net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_009 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M15 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M16 VDD RN net_003 VDD P_ISO W=0.475e-06 L=0.18e-06
M17 VDD D net_003 VDD P_ISO W=0.72e-06 L=0.18e-06
M18 net_004 net_001 net_003 VDD P_ISO W=0.41e-06 L=0.18e-06
M19 net_004 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 VDD net_006 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD net_004 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 net_007 net_000 net_006 VDD P_ISO W=0.6e-06 L=0.18e-06
M23 net_007 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M24 VDD net_009 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_007 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_009 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFFTR_X4_18_SVT_WB D RN CK Q QN VDD VSS
*.PININFO D:I RN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.66e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 VSS RN net_002 VSS N_ISO W=0.54e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.54e-06 L=0.18e-06
M4 net_004 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M5 net_004 net_001 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_006 net_005 VSS N_ISO W=0.22e-06 L=0.18e-06
M7 VSS net_004 net_006 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_007 net_001 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_007 net_000 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_007 net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_009 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_009 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 VDD net_000 net_001 VDD P_ISO W=0.75e-06 L=0.18e-06
M18 VDD RN net_003 VDD P_ISO W=0.475e-06 L=0.18e-06
M19 VDD D net_003 VDD P_ISO W=0.72e-06 L=0.18e-06
M20 net_004 net_001 net_003 VDD P_ISO W=0.41e-06 L=0.18e-06
M21 net_004 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_006 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M23 VDD net_004 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_007 net_000 net_006 VDD P_ISO W=0.615e-06 L=0.18e-06
M25 net_007 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_009 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_007 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD net_009 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_009 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DFF_X1_18_SVT_WB D CK Q QN VDD VSS
*.PININFO D:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.495e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.455e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M11 VSS net_006 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 VSS net_008 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M13 VDD CK net_000 VDD P_ISO W=0.48e-06 L=0.18e-06
M14 VDD net_000 net_001 VDD P_ISO W=0.65e-06 L=0.18e-06
M15 VDD net_001 net_009 VDD P_ISO W=0.605e-06 L=0.18e-06
M16 net_003 D net_009 VDD P_ISO W=0.605e-06 L=0.18e-06
M17 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M19 net_005 net_003 VDD VDD P_ISO W=0.47e-06 L=0.18e-06
M20 net_006 net_000 net_005 VDD P_ISO W=0.475e-06 L=0.18e-06
M21 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M23 VDD net_006 QN VDD P_ISO W=0.575e-06 L=0.18e-06
M24 VDD net_006 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_008 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DFF_X2_18_SVT_WB D CK Q QN VDD VSS
*.PININFO D:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.595e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.49e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.49e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.56e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.495e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 QN VSS N_ISO W=1.025e-06 L=0.18e-06
M11 VSS net_006 net_008 VSS N_ISO W=0.59e-06 L=0.18e-06
M12 VSS net_008 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M14 VDD net_000 net_001 VDD P_ISO W=0.945e-06 L=0.18e-06
M15 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M16 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M17 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M19 net_005 net_003 VDD VDD P_ISO W=0.665e-06 L=0.18e-06
M20 net_006 net_000 net_005 VDD P_ISO W=0.685e-06 L=0.18e-06
M21 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M23 VDD net_006 QN VDD P_ISO W=1.125e-06 L=0.18e-06
M24 VDD net_006 net_008 VDD P_ISO W=0.61e-06 L=0.18e-06
M25 VDD net_008 Q VDD P_ISO W=0.995e-06 L=0.18e-06
.ends

.subckt DFF_X4_18_SVT_WB D CK Q QN VDD VSS
*.PININFO D:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.595e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.49e-06 L=0.18e-06
M3 net_003 D net_002 VSS N_ISO W=0.49e-06 L=0.18e-06
M4 net_003 net_001 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.22e-06 L=0.18e-06
M6 VSS net_003 net_005 VSS N_ISO W=0.635e-06 L=0.18e-06
M7 net_006 net_001 net_005 VSS N_ISO W=0.545e-06 L=0.18e-06
M8 net_006 net_000 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 QN VSS N_ISO W=1.025e-06 L=0.18e-06
M11 VSS net_006 QN VSS N_ISO W=1.025e-06 L=0.18e-06
M12 VSS net_006 net_008 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_008 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_008 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VDD CK net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M16 VDD net_000 net_001 VDD P_ISO W=0.945e-06 L=0.18e-06
M17 VDD net_001 net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M18 net_003 D net_009 VDD P_ISO W=0.685e-06 L=0.18e-06
M19 net_003 net_000 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 VDD net_005 net_010 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 net_005 net_003 VDD VDD P_ISO W=0.685e-06 L=0.18e-06
M22 net_006 net_000 net_005 VDD P_ISO W=0.72e-06 L=0.18e-06
M23 net_006 net_001 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M24 VDD net_008 net_011 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_006 QN VDD P_ISO W=1.125e-06 L=0.18e-06
M26 VDD net_006 QN VDD P_ISO W=1.125e-06 L=0.18e-06
M27 VDD net_006 net_008 VDD P_ISO W=1.125e-06 L=0.18e-06
M28 VDD net_008 Q VDD P_ISO W=1.125e-06 L=0.18e-06
M29 VDD net_008 Q VDD P_ISO W=1.125e-06 L=0.18e-06
.ends

.subckt DLY1_X1_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.36e-06
M1 net_000 A net_001 VSS N_ISO W=0.42e-06 L=0.36e-06
M2 VSS net_001 Q VSS N_ISO W=0.52e-06 L=0.18e-06
M3 net_002 A net_001 VDD P_ISO W=0.42e-06 L=0.36e-06
M4 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.36e-06
M5 VDD net_001 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DLY1_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.36e-06
M1 net_000 A net_001 VSS N_ISO W=0.42e-06 L=0.36e-06
M2 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_002 A net_001 VDD P_ISO W=0.42e-06 L=0.36e-06
M5 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.36e-06
M6 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DLY2_X1_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.54e-06
M1 net_000 A net_001 VSS N_ISO W=0.42e-06 L=0.54e-06
M2 VSS net_001 Q VSS N_ISO W=0.52e-06 L=0.18e-06
M3 net_002 A net_001 VDD P_ISO W=0.42e-06 L=0.54e-06
M4 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.54e-06
M5 VDD net_001 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DLY2_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.54e-06
M1 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.54e-06
M2 Q net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_002 A net_001 VDD P_ISO W=0.42e-06 L=0.54e-06
M5 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.54e-06
M6 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DLY3_X1_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.72e-06
M1 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.72e-06
M2 VSS net_001 Q VSS N_ISO W=0.52e-06 L=0.18e-06
M3 net_001 A net_002 VDD P_ISO W=0.42e-06 L=0.72e-06
M4 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.72e-06
M5 VDD net_001 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DLY3_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.72e-06
M1 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.72e-06
M2 Q net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_001 A net_002 VDD P_ISO W=0.42e-06 L=0.72e-06
M5 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.72e-06
M6 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt DLY4_X1_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.9e-06
M1 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.9e-06
M2 VSS net_001 Q VSS N_ISO W=0.52e-06 L=0.18e-06
M3 net_001 A net_002 VDD P_ISO W=0.42e-06 L=0.9e-06
M4 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.9e-06
M5 VDD net_001 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt DLY4_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.32e-06 L=0.9e-06
M1 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.9e-06
M2 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_001 A net_002 VDD P_ISO W=0.42e-06 L=0.9e-06
M5 VDD A net_002 VDD P_ISO W=0.42e-06 L=0.9e-06
M6 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FA1_X0_18_SVT_WB A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
M0 VSS net_000 S VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_000 CI net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_004 net_003 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS A net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 net_004 B VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M7 VSS CI net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 VSS B net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_005 A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M10 net_003 CI net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 net_006 B net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 VSS A net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 CO net_003 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M14 VDD net_000 S VDD P_ISO W=0.42e-06 L=0.18e-06
M15 net_007 A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M16 net_008 B net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 net_000 CI net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 net_009 net_003 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD A net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 net_009 B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD CI net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD B net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 net_010 A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_003 CI net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 net_011 B net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD A net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 CO net_003 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt FA1_X1_18_SVT_WB A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
M0 VSS net_002 S VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_000 B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 CI net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_003 net_005 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS A net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS B net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_003 CI VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M8 VSS B net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 VSS A net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 net_005 CI net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 net_005 B net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 VSS A net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 VSS net_005 CO VSS N_ISO W=0.525e-06 L=0.18e-06
M14 VDD net_002 S VDD P_ISO W=0.575e-06 L=0.18e-06
M15 VDD A net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M16 net_007 B net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 net_002 CI net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 net_009 net_005 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD A net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD B net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 net_009 CI VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD B net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD A net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_005 CI net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 net_005 B net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD A net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD net_005 CO VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt FA1_X2_18_SVT_WB A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
M0 VSS net_002 S VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_000 B net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_002 CI net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 net_003 net_005 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS A net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS B net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M7 net_003 CI VSS VSS N_ISO W=0.44e-06 L=0.18e-06
M8 VSS B net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M9 VSS A net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M10 net_005 CI net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M11 net_005 B net_006 VSS N_ISO W=0.44e-06 L=0.18e-06
M12 VSS A net_006 VSS N_ISO W=0.44e-06 L=0.18e-06
M13 VSS net_005 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD net_002 S VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M16 net_007 B net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M17 net_002 CI net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M18 net_009 net_005 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M19 VDD A net_009 VDD P_ISO W=0.575e-06 L=0.18e-06
M20 VDD B net_009 VDD P_ISO W=0.575e-06 L=0.18e-06
M21 net_009 CI VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M22 VDD B net_010 VDD P_ISO W=0.575e-06 L=0.18e-06
M23 VDD A net_010 VDD P_ISO W=0.575e-06 L=0.18e-06
M24 net_005 CI net_010 VDD P_ISO W=0.575e-06 L=0.18e-06
M25 net_005 B net_011 VDD P_ISO W=0.575e-06 L=0.18e-06
M26 VDD A net_011 VDD P_ISO W=0.575e-06 L=0.18e-06
M27 VDD net_005 CO VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FA1_X4_18_SVT_WB A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
M0 VSS net_002 S VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_002 S VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_000 B net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 net_002 CI net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 net_003 net_005 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS A net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M7 VSS B net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M8 net_003 CI VSS VSS N_ISO W=0.44e-06 L=0.18e-06
M9 VSS B net_004 VSS N_ISO W=0.62e-06 L=0.18e-06
M10 VSS A net_004 VSS N_ISO W=0.535e-06 L=0.18e-06
M11 net_005 CI net_004 VSS N_ISO W=0.535e-06 L=0.18e-06
M12 net_005 B net_006 VSS N_ISO W=0.535e-06 L=0.18e-06
M13 VSS A net_006 VSS N_ISO W=0.535e-06 L=0.18e-06
M14 VSS net_005 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_005 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VDD net_002 S VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 S VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M19 net_007 B net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M20 net_002 CI net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M21 net_009 net_005 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M22 VDD A net_009 VDD P_ISO W=0.575e-06 L=0.18e-06
M23 VDD B net_009 VDD P_ISO W=0.575e-06 L=0.18e-06
M24 net_009 CI VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M25 VDD B net_010 VDD P_ISO W=1.02e-06 L=0.18e-06
M26 VDD A net_010 VDD P_ISO W=0.72e-06 L=0.18e-06
M27 net_005 CI net_010 VDD P_ISO W=0.72e-06 L=0.18e-06
M28 net_005 B net_011 VDD P_ISO W=0.72e-06 L=0.18e-06
M29 VDD A net_011 VDD P_ISO W=0.72e-06 L=0.18e-06
M30 VDD net_005 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_005 CO VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FA1_X8_18_SVT_WB A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VSS:B
M0 VSS net_002 S VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_002 S VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_002 S VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_002 S VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 net_000 B net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 net_002 CI net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M7 net_003 net_005 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M8 VSS A net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M9 VSS B net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M10 net_003 CI VSS VSS N_ISO W=0.44e-06 L=0.18e-06
M11 VSS B net_004 VSS N_ISO W=0.62e-06 L=0.18e-06
M12 VSS A net_004 VSS N_ISO W=0.535e-06 L=0.18e-06
M13 net_005 CI net_004 VSS N_ISO W=0.535e-06 L=0.18e-06
M14 net_005 B net_006 VSS N_ISO W=0.535e-06 L=0.18e-06
M15 VSS A net_006 VSS N_ISO W=0.535e-06 L=0.18e-06
M16 VSS net_005 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_005 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_005 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_005 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VDD net_002 S VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_002 S VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_002 S VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_002 S VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD A net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M25 net_007 B net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M26 net_002 CI net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M27 net_009 net_005 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M28 VDD A net_009 VDD P_ISO W=0.575e-06 L=0.18e-06
M29 VDD B net_009 VDD P_ISO W=0.575e-06 L=0.18e-06
M30 net_009 CI VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M31 VDD B net_010 VDD P_ISO W=1.02e-06 L=0.18e-06
M32 VDD A net_010 VDD P_ISO W=0.72e-06 L=0.18e-06
M33 net_005 CI net_010 VDD P_ISO W=0.72e-06 L=0.18e-06
M34 net_005 B net_011 VDD P_ISO W=0.72e-06 L=0.18e-06
M35 VDD A net_011 VDD P_ISO W=0.72e-06 L=0.18e-06
M36 VDD net_005 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_005 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD net_005 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_005 CO VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FILLCAP_X16_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
M0 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FILLCAP_X32_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
M0 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M26 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M30 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FILLCAP_X4_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
M0 net_000 net_003 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_003 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M3 net_003 net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FILLCAP_X64_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
M0 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M23 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M24 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M25 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M26 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M27 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M28 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M29 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M30 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M31 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M32 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M34 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M38 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M42 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M44 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M45 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M46 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M47 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M48 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M49 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M50 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M51 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M52 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M53 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M54 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M55 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M56 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M57 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M58 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M59 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M60 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M61 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M62 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M63 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FILLCAP_X8_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
M0 net_000 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_001 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt FILLER_X1_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
.ends

.subckt FILLER_X16_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
.ends

.subckt FILLER_X2_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
.ends

.subckt FILLER_X32_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
.ends

.subckt FILLER_X4_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
.ends

.subckt FILLER_X8_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
.ends

.subckt FILLTIE_18_SVT_WB VDD VSS
*.PININFO VDD:B VSS:B
.ends

.subckt HA1_X1_18_SVT_WB A B CO S VDD VSS
*.PININFO A:I B:I CO:O S:O VDD:B VSS:B
M0 VSS net_001 CO VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_001 B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_003 B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_002 A net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_001 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS net_003 S VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VDD net_001 CO VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD A net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_001 B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD B net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 net_003 A net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD net_001 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M13 VDD net_003 S VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt HA1_X2_18_SVT_WB A B CO S VDD VSS
*.PININFO A:I B:I CO:O S:O VDD:B VSS:B
M0 VSS net_001 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_003 B net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_002 A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_001 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VSS net_003 S VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD net_001 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_001 B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M10 VDD B net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_003 A net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD net_001 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD net_003 S VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt HA1_X4_18_SVT_WB A B CO S VDD VSS
*.PININFO A:I B:I CO:O S:O VDD:B VSS:B
M0 VSS net_001 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_001 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_002 A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_003 S VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 S VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD net_001 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_001 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_003 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_003 S VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_003 S VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt HA1_X8_18_SVT_WB A B CO S VDD VSS
*.PININFO A:I B:I CO:O S:O VDD:B VSS:B
M0 VSS net_001 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_001 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_001 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 CO VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_003 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_002 A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_001 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 S VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_003 S VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 S VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 S VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD net_001 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_001 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_001 CO VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 net_003 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_001 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_003 S VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_003 S VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_003 S VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_003 S VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt HOLD_X1_18_SVT_WB Q VDD VSS
*.PININFO Q:B VDD:B VSS:B
M0 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS Q net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VDD net_000 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M3 VDD Q net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_AO22_X0_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q_neg B0 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_0 A0 Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS x1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q Q_neg VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VDD B1 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_2 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q_neg A0 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_2 x1 Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD A1N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 Q Q_neg VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_AO22_X1_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q_neg B0 net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_0 A0 Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS x1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VDD B1 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_2 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q_neg A0 net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_2 x1 Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD A1N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_AO22_X2_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q_neg B0 net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_0 A0 Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS x1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD B1 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_2 B0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q_neg A0 net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_2 x1 Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M10 VDD A1N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_AO22_X4_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_1 B1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q_neg B0 net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0 A0 Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS x1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A1N x1 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD B1 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_2 B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q_neg A0 net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_2 x1 Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A1N x1 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_AOI21_X0_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q B0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_0 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS x1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A1N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q A0 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_1 x1 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_AOI21_X1_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q B0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_0 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS x1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A1N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 B0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q A0 net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_1 x1 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_AOI21_X2_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N x1 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS x1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A1N x1 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_1 B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q A0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_1 x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_AOI21_X4_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.515e-06 L=0.18e-06
M1 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_001 A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_001 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_001 net_003 VDD P_ISO W=0.81e-06 L=0.18e-06
M12 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_AOI21_X8_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.715e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 VDD B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_001 A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_001 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_001 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 net_003 VDD P_ISO W=0.815e-06 L=0.18e-06
M16 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_INV_B_OAI22_X0_18_SVT_WB A0 A1N B0 B1N Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1N:I Q:O VDD:B VSS:B
M0 VSS A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_001 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B1N net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q A1N net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VDD A0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B0 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD net_001 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q B1N net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 Q A1N net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD net_000 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_INV_B_OAI22_X1_18_SVT_WB A0 A1N B0 B1N Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1N:I Q:O VDD:B VSS:B
M0 VSS A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_001 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B1N net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_002 A1N Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 Q net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VDD A0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B0 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD net_001 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q B1N net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_004 A1N Q VDD P_ISO W=0.575e-06 L=0.18e-06
M11 VDD net_000 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_INV_B_OAI22_X2_18_SVT_WB A0 A1N B0 B1N Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1N:I Q:O VDD:B VSS:B
M0 VSS A0 x1 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 x2 B0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS x2 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 B1N VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A1N net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_0 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A0 x1 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 x2 B0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_2 x2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q B1N net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_1 A1N Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD x1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_INV_B_OAI22_X4_18_SVT_WB A0 A1N B0 B1N Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1N:I Q:O VDD:B VSS:B
M0 VSS B0 x2 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_0 x2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B1N net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 B1N VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS x2 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 x1 A0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q x1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_0 A1N Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A1N net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_0 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD B0 x2 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_2_0 x2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q B1N net_2_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_2_1 B1N Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD x2 net_2_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 x1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_1_0 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A1N net_1_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_1_1 A1N Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD x1 net_1_1 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND2_X0_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_NAND2_X1_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q net_000 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_NAND2_X12_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 x1 AN VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS AN x1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_0 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q x1 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_1 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_2 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q x1 net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_3 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B net_0_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_0_4 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q x1 net_0_4 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_0_5 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS B net_0_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 x1 AN VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD AN x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND2_X2_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD AN net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND2_X4_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD AN net_000 VDD P_ISO W=0.815e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND2_X8_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 x1 AN VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS AN x1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_0 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q x1 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_1 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_2 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q x1 net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_3 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B net_0_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 x1 AN VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD AN x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND3_X0_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_1 C VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_0 B net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q x1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD AN x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q C VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q x1 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_NAND3_X1_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_1 C VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_0 B net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q x1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD AN x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q C VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q x1 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_NAND3_X2_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS C net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD AN net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND3_X4_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN x1 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_1_0 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q x1 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_1 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_1_1 B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD AN x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND4_X0_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_2 D VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_1 C net_2 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_0 B net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q x1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD AN x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q D VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD C Q VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD x1 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_NAND4_X1_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_2 D VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_1 C net_2 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_0 B net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q x1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD AN x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q D VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD C Q VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD x1 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_NAND4_X2_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 C net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 B net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q net_000 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD AN net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NAND4_X4_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN x1 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_2_0 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_1_0 C net_2_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q x1 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_0_1 x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_1_1 B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_2_1 C net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS D net_2_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD AN x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD x1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR2_X0_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q net_000 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_NOR2_X1_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 Q net_000 net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_NOR2_X12_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_002 net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 Q net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_004 net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M25 Q net_000 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M26 net_006 net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD B net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR2_X2_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD AN net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M4 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR2_X4_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q net_000 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR2_X8_18_SVT_WB AN B Q VDD VSS
*.PININFO AN:I B:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_002 net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR3_X0_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD C net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_002 B net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q net_000 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_NOR3_X1_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD C net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_001 B net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q net_000 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_NOR3_X2_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD AN net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_002 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_002 net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR3_X4_18_SVT_WB AN B C Q VDD VSS
*.PININFO AN:I B:I C:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_002 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_003 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR4_X0_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS D Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q C VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD D net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_002 C net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_002 B net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q net_000 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_NOR4_X1_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS D Q VSS N_ISO W=0.575e-06 L=0.18e-06
M2 VSS C Q VSS N_ISO W=0.575e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.575e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=0.575e-06 L=0.18e-06
M5 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD D net_001 VDD P_ISO W=0.525e-06 L=0.18e-06
M7 net_002 C net_001 VDD P_ISO W=0.525e-06 L=0.18e-06
M8 net_003 B net_002 VDD P_ISO W=0.525e-06 L=0.18e-06
M9 net_003 net_000 Q VDD P_ISO W=0.525e-06 L=0.18e-06
.ends

.subckt INV_A_NOR4_X2_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD AN net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD D net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_002 C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_002 B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_NOR4_X4_18_SVT_WB AN B C D Q VDD VSS
*.PININFO AN:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD D net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_002 C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_002 B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_004 B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_006 C net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD D net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI211_X0_18_SVT_WB A0 A1N B0 C0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I C0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 C0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 B0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_002 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD C0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD net_000 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_OAI211_X1_18_SVT_WB A0 A1N B0 C0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I C0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS C0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 B0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_002 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD C0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q B0 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD net_000 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_OAI211_X2_18_SVT_WB A0 A1N B0 C0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I C0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS C0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI211_X4_18_SVT_WB A0 A1N B0 C0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I C0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS C0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_003 net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 A0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_003 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD C0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_003 A0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_003 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI21_X0_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q A0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_001 net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_OAI21_X1_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q A0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_001 net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD net_000 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_OAI21_X2_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_002 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI21_X4_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.475e-06 L=0.18e-06
M1 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_002 net_003 VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD A1N net_000 VDD P_ISO W=0.675e-06 L=0.18e-06
M8 VDD B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_004 A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_002 net_003 VDD P_ISO W=0.81e-06 L=0.18e-06
M12 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI21_X8_18_SVT_WB A0 A1N B0 Q VDD VSS
*.PININFO A0:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_002 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_002 net_003 VSS N_ISO W=0.715e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD A1N net_000 VDD P_ISO W=0.525e-06 L=0.18e-06
M11 VDD B0 net_002 VDD P_ISO W=1.05e-06 L=0.18e-06
M12 net_004 A0 net_002 VDD P_ISO W=1.05e-06 L=0.18e-06
M13 VDD net_000 net_004 VDD P_ISO W=1.05e-06 L=0.18e-06
M14 VDD net_002 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_002 net_003 VDD P_ISO W=0.815e-06 L=0.18e-06
M16 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI22_X0_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_001 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_001 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD net_000 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_A_OAI22_X1_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_001 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD net_000 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_A_OAI22_X2_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_001 net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_001 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI22_X4_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A1N net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_001 net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD A1N net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD B1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q B0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD B1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_A_OAI22_X8_18_SVT_WB A0 A1N B0 B1 Q VDD VSS
*.PININFO A0:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 net_002 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A1N net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A1N net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS A1N net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A1N net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_001 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_001 net_003 VSS N_ISO W=0.715e-06 L=0.18e-06
M10 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD B1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_001 B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_005 A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A1N net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD A1N net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD A1N net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD A1N net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_001 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_001 net_003 VDD P_ISO W=0.815e-06 L=0.18e-06
M24 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_B_AOI21_X0_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS B0N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q x1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_0 A1 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS A0 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD B0N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 x1 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q A1 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_1 A0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_B_AOI21_X1_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS B0N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q x1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_0 A1 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS A0 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD B0N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 x1 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q A1 net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_1 A0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_B_AOI21_X2_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS B0N x1 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q x1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A0 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD B0N x1 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_1 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q A1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_1 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_B_AOI21_X4_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 net_0 A0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 x1 A1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_1 x1 x2 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0N net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q x2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS x2 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 x1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A1 x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 x2 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B0N x2 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q x2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD x2 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_B_AOI21_X8_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 net_0 A0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 x1 A1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_1 x1 x2 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0N net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q x2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS x2 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q x2 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS x2 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 x1 A0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A1 x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 x2 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B0N x2 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q x2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD x2 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q x2 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD x2 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_B_OAI21_X0_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS B0N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 net_000 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q A1 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_001 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD B0N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q A1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_B_OAI21_X1_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS B0N net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 net_000 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q A1 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_001 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD B0N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q A1 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_B_OAI21_X2_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS B0N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD B0N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_B_OAI21_X4_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0N net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_000 A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_001 net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B0N net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_B_OAI21_X8_18_SVT_WB A0 A1 B0N Q VDD VSS
*.PININFO A0:I A1:I B0N:I Q:O VDD:B VSS:B
M0 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0N net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_000 A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_001 net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B0N net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X1_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X10_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=0.81e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.49e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.49e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.49e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.49e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.49e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.49e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X12_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.685e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.51e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.51e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.51e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.175e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.495e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.51e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.51e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=0.81e-06 L=0.18e-06
.ends

.subckt INVP2_X14_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.45e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.45e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.45e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.11e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.45e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.45e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.45e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.45e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=0.81e-06 L=0.18e-06
.ends

.subckt INVP2_X16_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M5 Q A VSS VSS N_ISO W=0.67e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=0.67e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M19 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M20 VDD A Q VDD P_ISO W=1.52e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X2_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X20_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M7 Q A VSS VSS N_ISO W=0.675e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M12 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M14 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M19 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M20 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M22 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M23 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M24 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M26 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M27 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M28 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M29 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X24_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M9 Q A VSS VSS N_ISO W=0.675e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M12 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M14 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M15 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M16 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M17 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M18 VSS A Q VSS N_ISO W=0.675e-06 L=0.18e-06
M19 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M22 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M23 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M24 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M26 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M27 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M28 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M29 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M30 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M31 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M32 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M33 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M34 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M35 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M36 VDD A Q VDD P_ISO W=1.525e-06 L=0.18e-06
M37 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X3_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.785e-06 L=0.18e-06
M1 Q A VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X5_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.875e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.875e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.875e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=0.805e-06 L=0.18e-06
M4 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X6_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.75e-06 L=0.18e-06
M4 VDD A Q VDD P_ISO W=0.805e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=1.445e-06 L=0.18e-06
M6 VDD A Q VDD P_ISO W=1.445e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=1.445e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INVP2_X8_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 VSS A Q VSS N_ISO W=0.7e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.7e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.7e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.7e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.7e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=0.815e-06 L=0.18e-06
M6 VDD A Q VDD P_ISO W=1.5e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=1.5e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.5e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.5e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=0.815e-06 L=0.18e-06
.ends

.subckt INV_X0_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt INV_X1_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt INV_X10_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A VDD VDD P_ISO W=0.805e-06 L=0.18e-06
M6 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X12_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=0.815e-06 L=0.18e-06
M8 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q A VDD VDD P_ISO W=0.815e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X14_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X16_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=0.81e-06 L=0.18e-06
M10 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X18_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M9 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A VDD VDD P_ISO W=0.81e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A VDD VDD P_ISO W=0.81e-06 L=0.18e-06
.ends

.subckt INV_X2_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X20_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.71e-06 L=0.18e-06
M10 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A VDD VDD P_ISO W=0.81e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD A Q VDD P_ISO W=0.81e-06 L=0.18e-06
.ends

.subckt INV_X24_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X3_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.785e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt INV_X32_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M15 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X4_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X5_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=0.875e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.875e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=0.875e-06 L=0.18e-06
M3 Q A VDD VDD P_ISO W=0.955e-06 L=0.18e-06
M4 VDD A Q VDD P_ISO W=0.955e-06 L=0.18e-06
M5 Q A VDD VDD P_ISO W=0.955e-06 L=0.18e-06
.ends

.subckt INV_X6_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt INV_X8_18_SVT_WB A Q VDD VSS
*.PININFO A:I Q:O VDD:B VSS:B
M0 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUX2_X0_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_003 net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q net_002 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_004 B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_002 net_000 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_005 S0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD A net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 Q net_002 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt MUX2_X1_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_003 net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q net_002 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_004 B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_002 net_000 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_005 S0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD A net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 Q net_002 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt MUX2_X12_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_002 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_005 S0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUX2_X2_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_003 net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 Q net_002 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_004 B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_002 net_000 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_005 S0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 VDD A net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 Q net_002 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUX2_X3_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_003 A VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=0.79e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=0.79e-06 L=0.18e-06
M7 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD B net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_002 net_000 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_002 S0 net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 VDD A net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=0.865e-06 L=0.18e-06
M13 VDD net_002 Q VDD P_ISO W=0.865e-06 L=0.18e-06
.ends

.subckt MUX2_X4_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD B net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_002 net_000 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_002 S0 net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 VDD A net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUX2_X6_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_002 net_000 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_002 S0 net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD A net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUX2_X8_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_002 net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_002 S0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_005 A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2D_X0_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 S0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_003 net_000 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q B net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_004 A Q VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD S0 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt MUXI2D_X1_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q A net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD net_000 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q B net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q A net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD S0 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt MUXI2D_X1P5_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M1 VSS S0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 B Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.555e-06 L=0.18e-06
M6 VDD S0 net_003 VDD P_ISO W=1.115e-06 L=0.18e-06
M7 Q A net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD net_000 net_004 VDD P_ISO W=1.115e-06 L=0.18e-06
.ends

.subckt MUXI2D_X2_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_001 S0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_003 net_000 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_004 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD S0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2D_X4_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS net_000 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD net_000 net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_002 B net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_002 A net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD S0 net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2D_X8_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS S0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_004 net_002 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD net_000 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_002 B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_006 A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD S0 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2PG_X4_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=0.9e-06 L=0.18e-06
M4 VSS S0 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q S0 net_001 VSS N_ISO W=0.9e-06 L=0.18e-06
M6 net_000 net_002 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M7 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD S0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 net_000 S0 Q VDD P_ISO W=1.3e-06 L=0.18e-06
M13 Q net_002 net_001 VDD P_ISO W=1.3e-06 L=0.18e-06
.ends

.subckt MUXI2PG_X6_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=0.88e-06 L=0.18e-06
M3 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M4 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M5 Q S0 net_001 VSS N_ISO W=0.88e-06 L=0.18e-06
M6 net_001 S0 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M7 VSS S0 net_002 VSS N_ISO W=0.88e-06 L=0.18e-06
M8 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M15 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M16 Q S0 net_000 VDD P_ISO W=1.32e-06 L=0.18e-06
M17 net_000 S0 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M18 VDD S0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2PG_X8_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A net_000 VSS N_ISO W=0.88e-06 L=0.18e-06
M4 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M5 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M6 Q S0 net_001 VSS N_ISO W=0.88e-06 L=0.18e-06
M7 net_001 S0 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M8 VSS S0 net_002 VSS N_ISO W=0.88e-06 L=0.18e-06
M9 VSS B net_001 VSS N_ISO W=0.88e-06 L=0.18e-06
M10 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M18 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M19 Q S0 net_000 VDD P_ISO W=1.32e-06 L=0.18e-06
M20 Q S0 net_000 VDD P_ISO W=1.32e-06 L=0.18e-06
M21 VDD S0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2_X0_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q S0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_003 B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q net_000 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_004 S0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD A net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt MUXI2_X1_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.555e-06 L=0.18e-06
M6 net_003 B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q net_000 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_004 S0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD A net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt MUXI2_X12_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M14 VDD B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_002 net_000 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_006 S0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2_X1P5_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 S0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.555e-06 L=0.18e-06
M6 VDD B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_003 net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_004 S0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2_X2_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_001 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q S0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_003 B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_004 S0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2_X3_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.785e-06 L=0.18e-06
M6 VSS net_004 Q VSS N_ISO W=0.785e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=0.785e-06 L=0.18e-06
M8 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_002 net_000 net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_006 S0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 net_006 A VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD net_002 net_004 VDD P_ISO W=0.865e-06 L=0.18e-06
M14 VDD net_004 Q VDD P_ISO W=0.865e-06 L=0.18e-06
M15 VDD net_004 Q VDD P_ISO W=0.865e-06 L=0.18e-06
.ends

.subckt MUXI2_X4_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_002 net_000 net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_006 S0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD A net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2_X6_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 S0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD S0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD B net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_002 net_000 net_005 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 net_006 S0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD A net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M14 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt MUXI2_X8_18_SVT_WB A B S0 Q VDD VSS
*.PININFO A:I B:I S0:I Q:O VDD:B VSS:B
M0 VSS S0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 S0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_002 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD S0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_002 net_000 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_006 S0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_A_NAND2_X0_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A0N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD net_000 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND2_A_NAND2_X1_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A0N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND2_A_NAND2_X2_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A0N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_A_NAND2_X4_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 net_001 A0N net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q B0 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A0N net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A1N net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_A_NOR3_X0_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 BN net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS AN net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS C Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS D Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD BN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD AN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_003 C net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_003 D Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND2_A_NOR3_X1_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 BN net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS AN net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS C Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS D Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD BN net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_000 AN VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_003 C net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q D net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND2_A_NOR3_X2_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 BN net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS AN net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD BN net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_000 AN VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_003 C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_003 D Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_A_NOR3_X4_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 BN net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS AN net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD BN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD AN net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_002 C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_004 D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_004 C net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_000 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_A_OAI21_X0_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 net_000 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_002 B1 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD A0N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD A1N net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND2_A_OAI21_X1_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 net_000 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_002 B1 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD A0N net_000 VDD P_ISO W=0.47e-06 L=0.18e-06
M6 VDD A1N net_000 VDD P_ISO W=0.47e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND2_A_OAI21_X2_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q B1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD A0N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD A1N net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_A_OAI21_X4_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_002 B1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q B1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_002 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A0N net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A1N net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_A_OAI21_X8_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 A0N net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A1N net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_003 B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 B1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_003 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_003 net_004 VSS N_ISO W=0.715e-06 L=0.18e-06
M7 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD A0N net_000 VDD P_ISO W=0.57e-06 L=0.18e-06
M12 VDD A1N net_000 VDD P_ISO W=0.57e-06 L=0.18e-06
M13 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_003 B0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_004 net_003 VDD VDD P_ISO W=1.05e-06 L=0.18e-06
M17 VDD net_003 net_004 VDD P_ISO W=0.715e-06 L=0.18e-06
M18 VDD net_004 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M19 VDD net_004 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M20 VDD net_004 Q VDD P_ISO W=1.05e-06 L=0.18e-06
M21 VDD net_004 Q VDD P_ISO W=1.05e-06 L=0.18e-06
.ends

.subckt NAND2T_X0_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 B VSS VSS N_ISO W=0.84e-06 L=0.18e-06
M1 net_000 A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VDD B Q VDD P_ISO W=0.42e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND2T_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VDD B Q VDD P_ISO W=0.575e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND2T_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.195e-06 L=0.18e-06
M2 VSS B net_000 VSS N_ISO W=1.195e-06 L=0.18e-06
M3 VSS B net_000 VSS N_ISO W=1.195e-06 L=0.18e-06
M4 VSS B net_000 VSS N_ISO W=1.195e-06 L=0.18e-06
M5 VSS B net_000 VSS N_ISO W=1.195e-06 L=0.18e-06
M6 VSS B net_000 VSS N_ISO W=1.195e-06 L=0.18e-06
M7 VSS B net_000 VSS N_ISO W=1.195e-06 L=0.18e-06
M8 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M15 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M17 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M18 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M20 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M21 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M22 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M23 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M24 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M25 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M26 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2T_X16_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M2 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M3 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M4 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M5 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M6 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M7 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M8 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M9 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M10 VSS B net_000 VSS N_ISO W=1.365e-06 L=0.18e-06
M11 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M18 net_001 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M22 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M23 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M24 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M25 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M26 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M27 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M28 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M29 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M30 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M31 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M32 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M33 VDD B Q VDD P_ISO W=0.7e-06 L=0.18e-06
M34 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2T_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2T_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2T_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.325e-06 L=0.18e-06
M2 VSS B net_000 VSS N_ISO W=1.325e-06 L=0.18e-06
M3 VSS B net_000 VSS N_ISO W=1.325e-06 L=0.18e-06
M4 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M9 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M10 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M11 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M12 Q B VDD VDD P_ISO W=0.69e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2T_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_000 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_X0_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VDD B Q VDD P_ISO W=0.42e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND2_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_000 A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VDD B Q VDD P_ISO W=0.575e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND2_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_0_0 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_1 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_2 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_3 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B net_0_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_4 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q A net_0_4 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_0_5 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B net_0_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_X16_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_0_0 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_0_1 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0_2 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_3 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B net_0_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_4 B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q A net_0_4 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_0_5 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B net_0_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_0_5 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS B net_0_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_0_5 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS B net_0_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M3 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_X24_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_004 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS B net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 Q A net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_007 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS B net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS B net_008 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 Q A net_008 VSS N_ISO W=1.05e-06 L=0.18e-06
M18 Q A net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS B net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS B net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M21 net_010 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M22 Q A net_011 VSS N_ISO W=1.05e-06 L=0.18e-06
M23 VSS B net_011 VSS N_ISO W=1.05e-06 L=0.18e-06
M24 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M42 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M44 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M45 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M46 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M47 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_X3_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_0_0 B VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M1 Q A net_0_0 VSS N_ISO W=0.785e-06 L=0.18e-06
M2 net_0_1 A Q VSS N_ISO W=0.785e-06 L=0.18e-06
M3 VSS B net_0_1 VSS N_ISO W=0.785e-06 L=0.18e-06
M4 Q B VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=0.86e-06 L=0.18e-06
M6 Q A VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M7 VDD B Q VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt NAND2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_X5_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 B VSS VSS N_ISO W=0.875e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=0.875e-06 L=0.18e-06
M2 net_001 A Q VSS N_ISO W=0.875e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=0.875e-06 L=0.18e-06
M4 net_002 B VSS VSS N_ISO W=0.875e-06 L=0.18e-06
M5 net_002 A Q VSS N_ISO W=0.875e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=0.955e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=0.955e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=0.955e-06 L=0.18e-06
M9 VDD B Q VDD P_ISO W=0.955e-06 L=0.18e-06
M10 VDD B Q VDD P_ISO W=0.955e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=0.955e-06 L=0.18e-06
.ends

.subckt NAND2_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3T_X0_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=0.84e-06 L=0.18e-06
M1 net_001 B net_000 VSS N_ISO W=0.84e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD C Q VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND3T_X1_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VDD C Q VDD P_ISO W=0.575e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND3T_X12_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_001 VSS N_ISO W=1.3e-06 L=0.18e-06
M2 VSS C net_002 VSS N_ISO W=1.3e-06 L=0.18e-06
M3 net_000 B net_002 VSS N_ISO W=1.3e-06 L=0.18e-06
M4 net_003 B net_000 VSS N_ISO W=1.3e-06 L=0.18e-06
M5 VSS C net_003 VSS N_ISO W=1.3e-06 L=0.18e-06
M6 VSS C net_004 VSS N_ISO W=1.3e-06 L=0.18e-06
M7 net_000 B net_004 VSS N_ISO W=1.3e-06 L=0.18e-06
M8 net_005 B net_000 VSS N_ISO W=1.3e-06 L=0.18e-06
M9 VSS C net_005 VSS N_ISO W=1.3e-06 L=0.18e-06
M10 VSS C net_006 VSS N_ISO W=1.3e-06 L=0.18e-06
M11 net_000 B net_006 VSS N_ISO W=1.3e-06 L=0.18e-06
M12 net_000 B net_007 VSS N_ISO W=1.3e-06 L=0.18e-06
M13 VSS C net_007 VSS N_ISO W=1.3e-06 L=0.18e-06
M14 VSS C net_008 VSS N_ISO W=1.3e-06 L=0.18e-06
M15 net_000 B net_008 VSS N_ISO W=1.3e-06 L=0.18e-06
M16 net_000 B net_009 VSS N_ISO W=1.3e-06 L=0.18e-06
M17 VSS C net_009 VSS N_ISO W=1.3e-06 L=0.18e-06
M18 VSS C net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M19 net_000 B net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M21 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M22 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M23 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M24 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M25 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M26 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M27 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M28 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M29 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M30 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M31 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M32 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M33 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M34 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M35 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M36 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M37 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M38 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M39 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M40 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M41 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M42 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M43 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M44 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M45 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M46 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M47 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M48 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M49 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M50 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3T_X16_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_001 VSS N_ISO W=1.27e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=1.27e-06 L=0.18e-06
M3 net_000 B net_002 VSS N_ISO W=1.27e-06 L=0.18e-06
M4 VSS C net_000 VSS N_ISO W=1.27e-06 L=0.18e-06
M5 VSS C net_003 VSS N_ISO W=1.27e-06 L=0.18e-06
M6 net_002 B net_003 VSS N_ISO W=1.27e-06 L=0.18e-06
M7 net_004 B net_002 VSS N_ISO W=1.27e-06 L=0.18e-06
M8 VSS C net_004 VSS N_ISO W=1.27e-06 L=0.18e-06
M9 VSS C net_005 VSS N_ISO W=1.27e-06 L=0.18e-06
M10 net_002 B net_005 VSS N_ISO W=1.27e-06 L=0.18e-06
M11 net_006 B net_002 VSS N_ISO W=1.27e-06 L=0.18e-06
M12 VSS C net_006 VSS N_ISO W=1.27e-06 L=0.18e-06
M13 VSS C net_007 VSS N_ISO W=1.27e-06 L=0.18e-06
M14 net_002 B net_007 VSS N_ISO W=1.27e-06 L=0.18e-06
M15 net_008 B net_002 VSS N_ISO W=1.27e-06 L=0.18e-06
M16 VSS C net_008 VSS N_ISO W=1.27e-06 L=0.18e-06
M17 VSS C net_009 VSS N_ISO W=1.27e-06 L=0.18e-06
M18 net_002 B net_009 VSS N_ISO W=1.27e-06 L=0.18e-06
M19 net_002 B net_010 VSS N_ISO W=1.27e-06 L=0.18e-06
M20 VSS C net_010 VSS N_ISO W=1.27e-06 L=0.18e-06
M21 VSS C net_011 VSS N_ISO W=1.27e-06 L=0.18e-06
M22 net_002 B net_011 VSS N_ISO W=1.27e-06 L=0.18e-06
M23 net_002 B net_012 VSS N_ISO W=1.27e-06 L=0.18e-06
M24 VSS C net_012 VSS N_ISO W=1.27e-06 L=0.18e-06
M25 VSS C net_013 VSS N_ISO W=1.05e-06 L=0.18e-06
M26 net_002 B net_013 VSS N_ISO W=1.05e-06 L=0.18e-06
M27 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M28 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M29 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M30 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M31 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M32 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M33 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M34 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M35 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M36 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M37 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M38 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M39 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M40 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M41 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M42 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M43 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M44 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M45 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M46 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M47 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M48 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M49 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M50 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M51 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M52 Q C VDD VDD P_ISO W=0.685e-06 L=0.18e-06
M53 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M54 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M55 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M56 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M57 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M58 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M59 VDD C Q VDD P_ISO W=0.685e-06 L=0.18e-06
M60 VDD B Q VDD P_ISO W=0.685e-06 L=0.18e-06
M61 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M62 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M63 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M64 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M65 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M66 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M67 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M68 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3T_X2_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_000 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_000 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3T_X4_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_000 VSS N_ISO W=1.26e-06 L=0.18e-06
M2 net_001 B net_000 VSS N_ISO W=1.26e-06 L=0.18e-06
M3 net_001 B net_002 VSS N_ISO W=1.26e-06 L=0.18e-06
M4 VSS C net_002 VSS N_ISO W=1.26e-06 L=0.18e-06
M5 VSS C net_003 VSS N_ISO W=1.26e-06 L=0.18e-06
M6 net_003 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD C Q VDD P_ISO W=0.77e-06 L=0.18e-06
M10 VDD B Q VDD P_ISO W=0.77e-06 L=0.18e-06
M11 VDD B Q VDD P_ISO W=0.77e-06 L=0.18e-06
M12 VDD C Q VDD P_ISO W=0.77e-06 L=0.18e-06
M13 VDD C Q VDD P_ISO W=0.77e-06 L=0.18e-06
M14 VDD B Q VDD P_ISO W=0.77e-06 L=0.18e-06
M15 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3T_X6_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_000 VSS N_ISO W=1.35e-06 L=0.18e-06
M2 VSS C net_000 VSS N_ISO W=1.35e-06 L=0.18e-06
M3 VSS C net_000 VSS N_ISO W=1.35e-06 L=0.18e-06
M4 VSS C net_000 VSS N_ISO W=1.35e-06 L=0.18e-06
M5 net_001 B net_000 VSS N_ISO W=1.35e-06 L=0.18e-06
M6 net_000 B net_001 VSS N_ISO W=1.35e-06 L=0.18e-06
M7 net_001 B net_000 VSS N_ISO W=1.35e-06 L=0.18e-06
M8 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_001 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_001 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M14 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M15 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M16 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M17 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M18 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M19 Q B VDD VDD P_ISO W=0.69e-06 L=0.18e-06
M20 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M21 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M22 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M23 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3T_X8_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 B net_000 VSS N_ISO W=1.37e-06 L=0.18e-06
M2 VSS C net_000 VSS N_ISO W=1.37e-06 L=0.18e-06
M3 VSS C net_002 VSS N_ISO W=1.37e-06 L=0.18e-06
M4 net_001 B net_002 VSS N_ISO W=1.37e-06 L=0.18e-06
M5 net_001 B net_003 VSS N_ISO W=1.37e-06 L=0.18e-06
M6 VSS C net_003 VSS N_ISO W=1.37e-06 L=0.18e-06
M7 VSS C net_004 VSS N_ISO W=1.37e-06 L=0.18e-06
M8 net_001 B net_004 VSS N_ISO W=1.37e-06 L=0.18e-06
M9 net_001 B net_005 VSS N_ISO W=1.37e-06 L=0.18e-06
M10 VSS C net_005 VSS N_ISO W=1.37e-06 L=0.18e-06
M11 VSS C net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_001 B net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 net_001 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M15 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VDD B Q VDD P_ISO W=0.765e-06 L=0.18e-06
M18 VDD B Q VDD P_ISO W=0.765e-06 L=0.18e-06
M19 VDD C Q VDD P_ISO W=0.765e-06 L=0.18e-06
M20 VDD C Q VDD P_ISO W=0.765e-06 L=0.18e-06
M21 VDD B Q VDD P_ISO W=0.765e-06 L=0.18e-06
M22 VDD C Q VDD P_ISO W=0.765e-06 L=0.18e-06
M23 VDD C Q VDD P_ISO W=0.765e-06 L=0.18e-06
M24 VDD B Q VDD P_ISO W=0.765e-06 L=0.18e-06
M25 VDD B Q VDD P_ISO W=0.765e-06 L=0.18e-06
M26 VDD C Q VDD P_ISO W=0.765e-06 L=0.18e-06
M27 VDD C Q VDD P_ISO W=0.765e-06 L=0.18e-06
M28 VDD B Q VDD P_ISO W=0.765e-06 L=0.18e-06
M29 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3_X0_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD C Q VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND3_X1_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_001 B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VDD C Q VDD P_ISO W=0.575e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND3_X12_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_1_5 B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_1_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_1_4 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 B net_1_4 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_1_3 B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_1_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_1_2 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_0 B net_1_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_1_1 B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS C net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_1_0 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_0_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 net_0 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 Q A net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M15 net_0 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 Q A net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 net_0 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3_X16_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_000 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 B net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 B net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_005 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS C net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS C net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_000 B net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_000 B net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS C net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS C net_008 VSS N_ISO W=1.05e-06 L=0.18e-06
M15 net_008 B net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 Q A net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M19 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M20 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M21 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M22 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M23 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M24 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M42 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M44 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M45 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M46 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M47 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3_X2_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_000 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3_X24_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_001 B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_000 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 B net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 B net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_000 B net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS C net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_006 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_000 B net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_000 B net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS C net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS C net_008 VSS N_ISO W=1.05e-06 L=0.18e-06
M15 net_000 B net_008 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 net_000 B net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS C net_009 VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS C net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M19 net_011 B net_010 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 Q A net_011 VSS N_ISO W=1.05e-06 L=0.18e-06
M21 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M22 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M23 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M24 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M25 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M26 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M27 net_000 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M28 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M29 Q A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M30 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M42 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M44 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M45 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M46 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M47 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M48 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M49 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M50 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M51 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M52 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M53 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M54 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M55 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M56 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M57 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M58 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M59 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3_X3_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_1_0 C VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M1 net_0_0 B net_1_0 VSS N_ISO W=0.785e-06 L=0.18e-06
M2 Q A net_0_0 VSS N_ISO W=0.785e-06 L=0.18e-06
M3 net_0_1 A Q VSS N_ISO W=0.785e-06 L=0.18e-06
M4 net_1_1 B net_0_1 VSS N_ISO W=0.785e-06 L=0.18e-06
M5 VSS C net_1_1 VSS N_ISO W=0.785e-06 L=0.18e-06
M6 Q C VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M7 VDD B Q VDD P_ISO W=0.86e-06 L=0.18e-06
M8 Q A VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=0.86e-06 L=0.18e-06
M10 Q B VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M11 VDD C Q VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt NAND3_X4_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_1_0 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_0_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0_1 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_1_1 B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3_X6_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_1_0 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_1_1 B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS C net_1_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_1_2 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_0_0 B net_1_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_0 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND3_X8_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 net_10 B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_10 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_11 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 B net_11 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_12 B net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_12 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_13 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_01 B net_13 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A net_01 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_0 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_0 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4T_X0_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 D VSS VSS N_ISO W=0.84e-06 L=0.18e-06
M1 net_001 C net_000 VSS N_ISO W=0.84e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=0.84e-06 L=0.18e-06
M3 Q A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q D VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD C Q VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q B VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND4T_X1_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q D VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD C Q VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q B VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND4T_X12_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M2 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M4 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M5 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M6 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M7 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M8 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M9 net_001 C net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M10 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M11 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M12 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M13 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M14 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M15 net_001 B net_002 VSS N_ISO W=1.455e-06 L=0.18e-06
M16 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M17 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M18 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M19 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M21 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M22 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M23 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M24 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M25 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M26 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M27 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M28 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M29 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M30 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M31 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M32 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M33 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M34 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M35 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M36 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M37 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M38 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M39 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M40 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M41 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M42 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M43 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M44 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M45 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M46 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M47 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M48 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M49 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M50 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M51 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M52 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M53 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4T_X16_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M2 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M4 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M5 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M6 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M7 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M8 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M9 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M10 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M11 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M12 VSS D net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M13 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M14 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M15 net_001 C net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M16 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M17 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M18 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M19 net_001 C net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M20 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M21 net_001 C net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M22 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M23 net_001 C net_000 VSS N_ISO W=1.455e-06 L=0.18e-06
M24 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M25 net_000 C net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M26 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M27 net_001 B net_002 VSS N_ISO W=1.455e-06 L=0.18e-06
M28 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M29 net_001 B net_002 VSS N_ISO W=1.455e-06 L=0.18e-06
M30 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M31 net_001 B net_002 VSS N_ISO W=1.455e-06 L=0.18e-06
M32 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M33 net_001 B net_002 VSS N_ISO W=1.455e-06 L=0.18e-06
M34 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M35 net_001 B net_002 VSS N_ISO W=1.455e-06 L=0.18e-06
M36 net_002 B net_001 VSS N_ISO W=1.455e-06 L=0.18e-06
M37 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M38 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M39 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M40 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M41 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M42 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M43 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M44 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M45 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M46 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M47 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M48 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M49 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M50 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M51 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M52 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M53 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M54 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M55 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M56 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M57 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M58 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M59 VDD D Q VDD P_ISO W=0.745e-06 L=0.18e-06
M60 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M61 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M62 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M63 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M64 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M65 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M66 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M67 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M68 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M69 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M70 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M71 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M72 VDD C Q VDD P_ISO W=0.745e-06 L=0.18e-06
M73 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M74 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M75 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M76 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M77 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M78 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M79 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M80 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M81 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M82 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M83 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M84 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M85 VDD B Q VDD P_ISO W=0.745e-06 L=0.18e-06
M86 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M87 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M88 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M89 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M90 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M91 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M92 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M93 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4T_X2_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_001_1 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000_1 C net_001_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS D net_000_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_000_0 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_001_0 C net_000_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_002 B net_001_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4T_X4_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_000 VSS N_ISO W=1.51e-06 L=0.18e-06
M2 VSS D net_000 VSS N_ISO W=1.51e-06 L=0.18e-06
M3 net_001 C net_000 VSS N_ISO W=1.51e-06 L=0.18e-06
M4 net_001 C net_000 VSS N_ISO W=1.51e-06 L=0.18e-06
M5 net_000 C net_001 VSS N_ISO W=1.51e-06 L=0.18e-06
M6 net_002 B net_001 VSS N_ISO W=1.51e-06 L=0.18e-06
M7 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M12 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M13 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M14 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M15 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M16 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M17 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M18 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M19 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M20 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4T_X6_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_000 VSS N_ISO W=1.315e-06 L=0.18e-06
M2 VSS D net_000 VSS N_ISO W=1.315e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=1.315e-06 L=0.18e-06
M4 VSS D net_000 VSS N_ISO W=1.315e-06 L=0.18e-06
M5 net_001 C net_000 VSS N_ISO W=1.315e-06 L=0.18e-06
M6 net_000 C net_001 VSS N_ISO W=1.315e-06 L=0.18e-06
M7 net_001 C net_000 VSS N_ISO W=1.315e-06 L=0.18e-06
M8 net_000 C net_001 VSS N_ISO W=1.315e-06 L=0.18e-06
M9 net_001 C net_000 VSS N_ISO W=1.315e-06 L=0.18e-06
M10 net_002 B net_001 VSS N_ISO W=1.315e-06 L=0.18e-06
M11 net_001 B net_002 VSS N_ISO W=1.315e-06 L=0.18e-06
M12 net_002 B net_001 VSS N_ISO W=1.315e-06 L=0.18e-06
M13 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M15 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M19 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M20 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M21 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M22 VDD D Q VDD P_ISO W=0.69e-06 L=0.18e-06
M23 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M24 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M25 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M26 VDD C Q VDD P_ISO W=0.69e-06 L=0.18e-06
M27 Q C VDD VDD P_ISO W=0.69e-06 L=0.18e-06
M28 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M29 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M30 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M31 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M32 VDD B Q VDD P_ISO W=0.69e-06 L=0.18e-06
M33 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4T_X8_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M2 VSS D net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M4 VSS D net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M5 VSS D net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M6 VSS D net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M7 net_001 C net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M8 net_000 C net_001 VSS N_ISO W=1.225e-06 L=0.18e-06
M9 net_001 C net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M10 net_000 C net_001 VSS N_ISO W=1.225e-06 L=0.18e-06
M11 net_001 C net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M12 net_000 C net_001 VSS N_ISO W=1.225e-06 L=0.18e-06
M13 net_001 C net_000 VSS N_ISO W=1.225e-06 L=0.18e-06
M14 net_002 B net_001 VSS N_ISO W=1.225e-06 L=0.18e-06
M15 net_001 B net_002 VSS N_ISO W=1.225e-06 L=0.18e-06
M16 net_002 B net_001 VSS N_ISO W=1.225e-06 L=0.18e-06
M17 net_001 B net_002 VSS N_ISO W=1.225e-06 L=0.18e-06
M18 net_002 B net_001 VSS N_ISO W=1.225e-06 L=0.18e-06
M19 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M21 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M22 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M23 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M24 Q A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M25 VDD D Q VDD P_ISO W=0.655e-06 L=0.18e-06
M26 VDD D Q VDD P_ISO W=0.655e-06 L=0.18e-06
M27 VDD D Q VDD P_ISO W=0.655e-06 L=0.18e-06
M28 VDD D Q VDD P_ISO W=0.655e-06 L=0.18e-06
M29 VDD D Q VDD P_ISO W=0.655e-06 L=0.18e-06
M30 VDD D Q VDD P_ISO W=0.655e-06 L=0.18e-06
M31 VDD D Q VDD P_ISO W=0.655e-06 L=0.18e-06
M32 VDD C Q VDD P_ISO W=0.655e-06 L=0.18e-06
M33 VDD C Q VDD P_ISO W=0.655e-06 L=0.18e-06
M34 VDD C Q VDD P_ISO W=0.655e-06 L=0.18e-06
M35 VDD C Q VDD P_ISO W=0.655e-06 L=0.18e-06
M36 VDD C Q VDD P_ISO W=0.655e-06 L=0.18e-06
M37 VDD C Q VDD P_ISO W=0.655e-06 L=0.18e-06
M38 VDD C Q VDD P_ISO W=0.655e-06 L=0.18e-06
M39 VDD B Q VDD P_ISO W=0.655e-06 L=0.18e-06
M40 VDD B Q VDD P_ISO W=0.655e-06 L=0.18e-06
M41 VDD B Q VDD P_ISO W=0.655e-06 L=0.18e-06
M42 VDD B Q VDD P_ISO W=0.655e-06 L=0.18e-06
M43 VDD B Q VDD P_ISO W=0.655e-06 L=0.18e-06
M44 VDD B Q VDD P_ISO W=0.655e-06 L=0.18e-06
M45 VDD B Q VDD P_ISO W=0.655e-06 L=0.18e-06
M46 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M47 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M48 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M49 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4_X0_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 C net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD D Q VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD C Q VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NAND4_X1_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_000 C net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q A net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD D Q VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD C Q VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NAND4_X12_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_2_0 C net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_2_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_2_1 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_1 C net_2_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_2_2 C net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS D net_2_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_2_3 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_1 C net_2_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_2_4 C net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS D net_2_4 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_2_5 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_1_0 C net_2_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_0_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_0_1 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 net_1 B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 net_0_2 B net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 Q A net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M18 net_0_3 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 net_1 B net_0_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M20 net_0_4 B net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M21 Q A net_0_4 VSS N_ISO W=1.05e-06 L=0.18e-06
M22 net_0_5 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M23 net_1 B net_0_5 VSS N_ISO W=1.05e-06 L=0.18e-06
M24 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M42 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M44 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M45 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M46 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M47 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4_X2_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_002 B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4_X4_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_000 C net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS D net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_003 C net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_004 B net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_004 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 B net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4_X6_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_2_0 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_1 C net_2_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_2_1 C net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS D net_2_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_2_2 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_1_0 C net_2_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_0_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_1 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_1 B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_0_2 B net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q A net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NAND4_X8_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 net_2_0 C net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D net_2_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_2_1 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_1 C net_2_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_2_2 C net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS D net_2_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_2_3 D VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_1_0 C net_2_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_0 B net_1_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q A net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_0_1 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_1 B net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_0_2 B net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 Q A net_0_2 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_0_3 A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 net_1 B net_0_3 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q D VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 Q B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M30 Q A VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M31 VDD B Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_AOI21_X0_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 x1 A0N VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_0 B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS B1 net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_2 A0N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD A1N net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_1 x1 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q B0 net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_1 B1 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NOR2_A_AOI21_X1_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 x1 A0N VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_0 B0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS B1 net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_2 A0N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD A1N net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_1 x1 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B0 net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 net_1 B1 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NOR2_A_AOI21_X2_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 x1 A0N VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A1N x1 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B1 net_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_2 A0N x1 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD A1N net_2 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_1 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_1 B1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_AOI21_X4_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 x1 A0N VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1N x1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0_1 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B1 net_0_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_0_0 B1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q B0 net_0_0 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_2 A0N x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A1N net_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_1 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q B0 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_1 B1 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q B1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_1 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD x1 net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_AOI21_X8_18_SVT_WB A0N A1N B0 B1 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A0N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A1N net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B1 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_003 net_001 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 net_003 VSS N_ISO W=0.715e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_000 A0N net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD A1N net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD net_000 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_001 B0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_001 B1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_001 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_001 net_003 VDD P_ISO W=0.815e-06 L=0.18e-06
M18 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_NAND3_X0_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 x1 BN VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS AN x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_1 x1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_0 C net_1 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q D net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_2 BN x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD AN net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q x1 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD C Q VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q D VDD VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NOR2_A_NAND3_X1_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 x1 BN VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS AN x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_1 x1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_0 C net_1 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q D net_0 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_2 BN x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD AN net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q x1 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD C Q VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q D VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NOR2_A_NAND3_X2_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 VSS BN net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_000 AN VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 C net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_002 D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 BN net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD AN net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_NAND3_X4_18_SVT_WB AN BN C D Q VDD VSS
*.PININFO AN:I BN:I C:I D:I Q:O VDD:B VSS:B
M0 VSS BN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS AN net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 C net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q D net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_003 D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_003 C net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_000 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_000 BN net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD AN net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD D Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD C Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_NOR2_X0_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 x1 A0N VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_1 A0N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD A1N net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_0 x1 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q B0 net_0 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NOR2_A_NOR2_X1_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 x1 A0N VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A1N x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_1 A0N x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD A1N net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_0 x1 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q B0 net_0 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NOR2_A_NOR2_X2_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 x1 A0N VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A1N x1 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_1 A0N x1 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD A1N net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_0 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q B0 net_0 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_NOR2_X4_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 VSS A0N net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1N net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_001 A0N net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A1N net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_002 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_A_NOR2_X8_18_SVT_WB A0N A1N B0 Q VDD VSS
*.PININFO A0N:I A1N:I B0:I Q:O VDD:B VSS:B
M0 x1 A1N VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A0N x1 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 x1 A0N VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1N x1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q x1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q x1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS x1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_1_0_0 A1N VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 x1 A0N net_1_0_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_1_0_1 A0N x1 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A1N net_1_0_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_0_0_0 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q B0 net_0_0_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_0_0_1 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD x1 net_0_0_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 net_0_0_2 x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 Q B0 net_0_0_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_0_0_3 B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD x1 net_0_0_3 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3T_X10_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M6 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M12 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M14 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M15 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M16 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M17 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M18 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M19 net_000 A Q VDD P_ISO W=1.65e-06 L=0.18e-06
M20 net_000 A Q VDD P_ISO W=1.65e-06 L=0.18e-06
M21 Q A net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M22 net_000 A Q VDD P_ISO W=1.65e-06 L=0.18e-06
M23 net_000 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3T_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.45e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.45e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.45e-06 L=0.18e-06
M3 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 VDD B net_000 VDD P_ISO W=1.55e-06 L=0.18e-06
M5 net_000 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3T_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.5e-06 L=0.18e-06
M1 Q B VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.5e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.5e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=0.5e-06 L=0.18e-06
M5 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B net_000 VDD P_ISO W=1.58e-06 L=0.18e-06
M7 VDD B net_000 VDD P_ISO W=1.58e-06 L=0.18e-06
M8 Q A net_000 VDD P_ISO W=1.58e-06 L=0.18e-06
M9 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3T_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q B VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.5e-06 L=0.18e-06
M2 Q B VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.5e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.5e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M7 VDD B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_005 B VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M9 VDD B net_005 VDD P_ISO W=1.66e-06 L=0.18e-06
M10 net_005 B VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M11 Q A net_005 VDD P_ISO W=1.66e-06 L=0.18e-06
M12 net_005 A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M13 Q A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.22e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VDD B net_000 VDD P_ISO W=0.66e-06 L=0.18e-06
M3 Q A net_000 VDD P_ISO W=0.66e-06 L=0.18e-06
.ends

.subckt NOR2P3_X14_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M6 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M12 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M14 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M16 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M17 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M18 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M19 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M20 VDD B net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M21 Q A net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M22 net_000 A Q VDD P_ISO W=1.65e-06 L=0.18e-06
M23 Q A net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M24 net_000 A Q VDD P_ISO W=1.65e-06 L=0.18e-06
M25 Q A net_000 VDD P_ISO W=1.65e-06 L=0.18e-06
M26 net_000 A Q VDD P_ISO W=1.65e-06 L=0.18e-06
M27 net_000 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3_X16_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M6 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M7 VSS B Q VSS N_ISO W=0.55e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M12 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M14 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M15 VSS A Q VSS N_ISO W=0.55e-06 L=0.18e-06
M16 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD B net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M18 VDD B net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M19 VDD B net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M20 VDD B net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M21 VDD B net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M22 VDD B net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M23 VDD B net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M24 Q A net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M25 net_000 A Q VDD P_ISO W=1.64e-06 L=0.18e-06
M26 Q A net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M27 net_000 A Q VDD P_ISO W=1.64e-06 L=0.18e-06
M28 Q A net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M29 net_000 A Q VDD P_ISO W=1.64e-06 L=0.18e-06
M30 Q A net_000 VDD P_ISO W=1.64e-06 L=0.18e-06
M31 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M3 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.45e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.45e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.45e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.45e-06 L=0.18e-06
M4 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD B net_000 VDD P_ISO W=1.55e-06 L=0.18e-06
M6 Q A net_000 VDD P_ISO W=1.55e-06 L=0.18e-06
M7 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q B VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.5e-06 L=0.18e-06
M2 Q B VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.5e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.5e-06 L=0.18e-06
M6 net_006 B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B net_006 VDD P_ISO W=1.66e-06 L=0.18e-06
M8 net_006 B VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M9 Q A net_006 VDD P_ISO W=1.66e-06 L=0.18e-06
M10 net_006 A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M11 Q A net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2P3_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q B VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.5e-06 L=0.18e-06
M2 Q B VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.5e-06 L=0.18e-06
M4 Q A VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.5e-06 L=0.18e-06
M6 Q A VSS VSS N_ISO W=0.5e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=0.5e-06 L=0.18e-06
M8 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_004 B VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M10 VDD B net_004 VDD P_ISO W=1.66e-06 L=0.18e-06
M11 net_004 B VDD VDD P_ISO W=1.66e-06 L=0.18e-06
M12 Q A net_004 VDD P_ISO W=1.66e-06 L=0.18e-06
M13 net_004 A Q VDD P_ISO W=1.66e-06 L=0.18e-06
M14 Q A net_004 VDD P_ISO W=1.66e-06 L=0.18e-06
M15 net_004 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_X0_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VDD B net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M3 net_000 A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NOR2_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VDD B net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M3 net_000 A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NOR2_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_001 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 Q A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M3 net_000 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_X3_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_X5_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=0.89e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=0.89e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.89e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=0.89e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=0.89e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=0.89e-06 L=0.18e-06
M6 VDD B net_000 VDD P_ISO W=0.955e-06 L=0.18e-06
M7 Q A net_000 VDD P_ISO W=0.955e-06 L=0.18e-06
M8 net_001 A Q VDD P_ISO W=0.955e-06 L=0.18e-06
M9 VDD B net_001 VDD P_ISO W=0.955e-06 L=0.18e-06
M10 VDD B net_002 VDD P_ISO W=0.955e-06 L=0.18e-06
M11 net_002 A Q VDD P_ISO W=0.955e-06 L=0.18e-06
.ends

.subckt NOR2_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_001 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR3_X0_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C Q VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD C net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M4 net_001 B net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_001 A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NOR3_X1_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C Q VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VDD C net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M4 net_001 B net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_001 A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NOR3_X12_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 net_000 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_000 B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_000 B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD C net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M25 net_000 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M26 net_000 B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD C net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD C net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M29 net_006 B net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M30 Q A net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M31 net_000 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M32 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M33 net_000 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M34 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M35 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR3_X2_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 net_000 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR3_X4_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_001 B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_001 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_003 B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR3_X6_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_001 B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_001 B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_003 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_001 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_001 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR3_X8_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_000 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_000 B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_000 B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD C net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_005 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_000 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 Q A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR4_X0_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D Q VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD D net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_001 C net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_002 B net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_002 A Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt NOR4_X1_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D Q VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD D net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_001 C net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_002 B net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_002 A Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt NOR4_X12_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M23 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M24 net_000 C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD D net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD D net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M27 net_000 C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M28 net_003 C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M30 VDD D net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M31 net_000 C net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M32 net_000 C net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD D net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD D net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M35 net_007 C net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M36 net_008 B net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M37 net_008 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M38 Q A net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M39 net_000 B net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M40 net_010 B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M41 Q A net_010 VDD P_ISO W=1.15e-06 L=0.18e-06
M42 net_011 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M43 net_000 B net_011 VDD P_ISO W=1.15e-06 L=0.18e-06
M44 net_000 B net_012 VDD P_ISO W=1.15e-06 L=0.18e-06
M45 Q A net_012 VDD P_ISO W=1.15e-06 L=0.18e-06
M46 Q A net_013 VDD P_ISO W=1.15e-06 L=0.18e-06
M47 net_000 B net_013 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR4_X2_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD D net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 net_001 C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_001 B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_002 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR4_X4_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD D net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_001 C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_002 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_004 B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_005 C net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD D net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR4_X6_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD D net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_001 C net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_001 C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD D net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_004 C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_005 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q A net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q A net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_001 B net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_007 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 net_007 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt NOR4_X8_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS D Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS C Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS A Q VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M16 net_000 C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD D net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD D net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_000 C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 net_000 C net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD D net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 net_005 C net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 net_005 B net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M25 net_006 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q A net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M27 net_000 B net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M28 net_000 B net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M29 Q A net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M30 Q A net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M31 net_000 B net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OA21_X0_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 A0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_001 B0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_000 A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B0 net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OA21_X1_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 A0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_001 B0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_000 A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_000 B0 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OA21_X2_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=0.51e-06 L=0.18e-06
M1 net_000 A0 net_001 VSS N_ISO W=0.51e-06 L=0.18e-06
M2 net_001 B0 VSS VSS N_ISO W=0.575e-06 L=0.18e-06
M3 VSS net_000 Q VSS N_ISO W=1.045e-06 L=0.18e-06
M4 VDD A1 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_000 A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OA21_X4_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_001 A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OA21_X8_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=0.51e-06 L=0.18e-06
M1 net_000 A0 net_001 VSS N_ISO W=0.51e-06 L=0.18e-06
M2 VSS B0 net_001 VSS N_ISO W=0.575e-06 L=0.18e-06
M3 VSS net_000 net_002 VSS N_ISO W=1.045e-06 L=0.18e-06
M4 VSS net_002 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_002 net_003 VSS N_ISO W=0.715e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD A1 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 net_000 A0 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 VDD B0 net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD net_000 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_002 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_002 net_003 VDD P_ISO W=0.815e-06 L=0.18e-06
M16 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OA22_X0_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS net_001 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_001 A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_000 A1 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD net_001 Q VDD P_ISO W=0.58e-06 L=0.18e-06
M6 VDD B1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_001 B0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_001 A0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD A1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OA22_X1_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=0.425e-06 L=0.18e-06
M1 net_001 A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VSS B1 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD A1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_000 A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_000 B0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OA22_X2_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_001 A0 net_000 VSS N_ISO W=0.45e-06 L=0.18e-06
M2 VSS B0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS B1 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD A1 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_000 A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_000 B0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OA22_X4_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_001 A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_001 A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_000 A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_000 B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OA22_X8_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_001 A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_001 A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_001 A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_001 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M12 VDD B1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_001 B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_001 B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_001 A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_001 A0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD A1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_001 Q VDD P_ISO W=0.81e-06 L=0.18e-06
.ends

.subckt OAI12P2_X0_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_000 A1 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_000 B0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD A1 net_001 VDD P_ISO W=0.84e-06 L=0.18e-06
M4 Q A0 net_001 VDD P_ISO W=0.84e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.84e-06 L=0.18e-06
.ends

.subckt OAI12P2_X1_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_000 A1 Q VSS N_ISO W=0.55e-06 L=0.18e-06
M1 Q A0 net_000 VSS N_ISO W=0.55e-06 L=0.18e-06
M2 net_000 B0 VSS VSS N_ISO W=0.55e-06 L=0.18e-06
M3 VDD A1 net_002 VDD P_ISO W=1.1e-06 L=0.18e-06
M4 Q A0 net_002 VDD P_ISO W=1.1e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=1.1e-06 L=0.18e-06
.ends

.subckt OAI12P2_X10_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M1 net_000 A1 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M2 Q A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M3 net_000 A1 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M4 Q A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M5 net_000 A0 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M6 Q A0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M7 net_000 A0 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M8 Q A0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M9 net_000 A0 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M10 VSS B0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M11 VSS B0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M12 VSS B0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M13 VSS B0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M14 VSS B0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M15 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A1 net_001 VDD P_ISO W=1.395e-06 L=0.18e-06
M17 VDD A1 net_001 VDD P_ISO W=1.395e-06 L=0.18e-06
M18 VDD A1 net_001 VDD P_ISO W=1.395e-06 L=0.18e-06
M19 VDD A1 net_001 VDD P_ISO W=1.395e-06 L=0.18e-06
M20 Q A0 net_001 VDD P_ISO W=1.395e-06 L=0.18e-06
M21 net_001 A0 Q VDD P_ISO W=1.395e-06 L=0.18e-06
M22 Q A0 net_001 VDD P_ISO W=1.395e-06 L=0.18e-06
M23 net_001 A0 Q VDD P_ISO W=1.395e-06 L=0.18e-06
M24 Q A0 net_001 VDD P_ISO W=1.395e-06 L=0.18e-06
M25 VDD B0 Q VDD P_ISO W=1.395e-06 L=0.18e-06
M26 VDD B0 Q VDD P_ISO W=1.395e-06 L=0.18e-06
M27 VDD B0 Q VDD P_ISO W=1.395e-06 L=0.18e-06
M28 VDD B0 Q VDD P_ISO W=1.395e-06 L=0.18e-06
M29 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI12P2_X14_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M1 net_000 A1 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M2 Q A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M3 net_000 A1 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M4 Q A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M5 net_000 A1 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M6 Q A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M7 net_000 A0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M8 Q A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M9 net_000 A0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M10 Q A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M11 net_000 A0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M12 Q A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M13 net_000 A0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M14 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M15 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M16 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M17 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M18 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M19 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M20 net_000 B0 VSS VSS N_ISO W=0.715e-06 L=0.18e-06
M21 net_001 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_001 A1 VDD VDD P_ISO W=1.38e-06 L=0.18e-06
M23 net_001 A1 VDD VDD P_ISO W=1.38e-06 L=0.18e-06
M24 VDD A1 net_001 VDD P_ISO W=1.38e-06 L=0.18e-06
M25 net_001 A1 VDD VDD P_ISO W=1.38e-06 L=0.18e-06
M26 VDD A1 net_001 VDD P_ISO W=1.38e-06 L=0.18e-06
M27 net_001 A1 VDD VDD P_ISO W=1.38e-06 L=0.18e-06
M28 Q A0 net_001 VDD P_ISO W=1.38e-06 L=0.18e-06
M29 net_001 A0 Q VDD P_ISO W=1.38e-06 L=0.18e-06
M30 Q A0 net_001 VDD P_ISO W=1.38e-06 L=0.18e-06
M31 net_001 A0 Q VDD P_ISO W=1.38e-06 L=0.18e-06
M32 Q A0 net_001 VDD P_ISO W=1.38e-06 L=0.18e-06
M33 net_001 A0 Q VDD P_ISO W=1.38e-06 L=0.18e-06
M34 Q A0 net_001 VDD P_ISO W=1.38e-06 L=0.18e-06
M35 VDD B0 Q VDD P_ISO W=1.38e-06 L=0.18e-06
M36 Q B0 VDD VDD P_ISO W=1.38e-06 L=0.18e-06
M37 VDD B0 Q VDD P_ISO W=1.38e-06 L=0.18e-06
M38 Q B0 VDD VDD P_ISO W=1.38e-06 L=0.18e-06
M39 VDD B0 Q VDD P_ISO W=1.38e-06 L=0.18e-06
M40 Q B0 VDD VDD P_ISO W=1.38e-06 L=0.18e-06
M41 Q B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI12P2_X6_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M1 net_000 A1 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M2 net_000 A1 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M3 net_000 A0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M4 Q A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M5 net_000 A0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M6 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M7 VSS B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M8 net_000 B0 VSS VSS N_ISO W=0.715e-06 L=0.18e-06
M9 net_001 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A1 net_001 VDD P_ISO W=1.425e-06 L=0.18e-06
M11 VDD A1 net_001 VDD P_ISO W=1.425e-06 L=0.18e-06
M12 Q A0 net_001 VDD P_ISO W=1.425e-06 L=0.18e-06
M13 net_001 A0 Q VDD P_ISO W=1.425e-06 L=0.18e-06
M14 Q A0 net_001 VDD P_ISO W=1.425e-06 L=0.18e-06
M15 VDD B0 Q VDD P_ISO W=1.425e-06 L=0.18e-06
M16 VDD B0 Q VDD P_ISO W=1.425e-06 L=0.18e-06
M17 Q B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI12_X0_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A1 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M4 Q A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI12_X1_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_000 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 A1 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M4 Q A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI12_X2_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M4 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI12_X3_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS B0 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M2 Q A1 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M3 net_000 A0 Q VSS N_ISO W=0.79e-06 L=0.18e-06
M4 Q A0 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M5 Q A1 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M6 VDD B0 Q VDD P_ISO W=0.865e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=0.865e-06 L=0.18e-06
M8 VDD A1 net_001 VDD P_ISO W=0.865e-06 L=0.18e-06
M9 Q A0 net_001 VDD P_ISO W=0.865e-06 L=0.18e-06
M10 Q A0 net_002 VDD P_ISO W=0.865e-06 L=0.18e-06
M11 VDD A1 net_002 VDD P_ISO W=0.865e-06 L=0.18e-06
.ends

.subckt OAI12_X4_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_000 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_001_0 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A0 net_001_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_001_1 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A1 net_001_1 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI12_X6_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_000 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_001 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI12_X8_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 net_000 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_000 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_000 B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_000 B0 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_001 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_002 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_003 A1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_004 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q B0 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI211_X0_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 net_000 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_000 B0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q C0 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q A0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD C0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI211_X1_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 net_000 A1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_000 B0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q C0 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD A1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 Q A0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD C0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI211_X2_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_000 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q C0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI211_X4_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q C0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q C0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 B0 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI211_X8_18_SVT_WB A0 A1 B0 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I C0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_000 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_002 C0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_002 net_003 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_002 net_003 VSS N_ISO W=0.715e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_002 A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_002 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_002 net_003 VDD P_ISO W=0.815e-06 L=0.18e-06
M16 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI21P2_X0_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_000 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_000 B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD A1 net_002 VDD P_ISO W=0.84e-06 L=0.18e-06
M4 Q A0 net_002 VDD P_ISO W=0.84e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.84e-06 L=0.18e-06
.ends

.subckt OAI21P2_X1_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_000 A1 VSS VSS N_ISO W=0.55e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=0.55e-06 L=0.18e-06
M2 net_000 B0 Q VSS N_ISO W=0.55e-06 L=0.18e-06
M3 VDD A1 net_002 VDD P_ISO W=1.1e-06 L=0.18e-06
M4 Q A0 net_002 VDD P_ISO W=1.1e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=1.1e-06 L=0.18e-06
.ends

.subckt OAI21P2_X10_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M2 VSS A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M3 VSS A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M4 VSS A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M5 net_000 A0 VSS VSS N_ISO W=0.71e-06 L=0.18e-06
M6 VSS A0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M7 VSS A0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M8 VSS A0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M9 VSS A0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M10 Q B0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M11 net_000 B0 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M12 Q B0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M13 net_000 B0 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M14 net_000 B0 Q VSS N_ISO W=0.71e-06 L=0.18e-06
M15 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A1 net_001 VDD P_ISO W=1.41e-06 L=0.18e-06
M17 VDD A1 net_001 VDD P_ISO W=1.41e-06 L=0.18e-06
M18 VDD A1 net_001 VDD P_ISO W=1.41e-06 L=0.18e-06
M19 VDD A1 net_001 VDD P_ISO W=1.41e-06 L=0.18e-06
M20 net_001 A0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M21 net_001 A0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M22 Q A0 net_001 VDD P_ISO W=1.41e-06 L=0.18e-06
M23 net_001 A0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M24 net_001 A0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M25 VDD B0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M26 VDD B0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M27 VDD B0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M28 VDD B0 Q VDD P_ISO W=1.41e-06 L=0.18e-06
M29 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI21P2_X14_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M2 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M3 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M4 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M5 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M6 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M7 net_000 A0 VSS VSS N_ISO W=0.715e-06 L=0.18e-06
M8 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M9 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M10 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M11 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M12 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M13 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M14 Q B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M15 net_000 B0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M16 Q B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M17 net_000 B0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M18 Q B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M19 net_000 B0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M20 net_000 B0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M21 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD A1 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M23 VDD A1 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M24 VDD A1 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M25 VDD A1 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M26 VDD A1 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M27 VDD A1 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M28 Q A0 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M29 net_001 A0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M30 net_001 A0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M31 net_001 A0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M32 Q A0 net_001 VDD P_ISO W=1.39e-06 L=0.18e-06
M33 net_001 A0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M34 net_001 A0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M35 VDD B0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M36 VDD B0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M37 VDD B0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M38 VDD B0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M39 VDD B0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M40 VDD B0 Q VDD P_ISO W=1.39e-06 L=0.18e-06
M41 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI21P2_X6_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M2 VSS A1 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M3 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M4 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M5 VSS A0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M6 Q B0 net_000 VSS N_ISO W=0.715e-06 L=0.18e-06
M7 net_000 B0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M8 net_000 B0 Q VSS N_ISO W=0.715e-06 L=0.18e-06
M9 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A1 net_001 VDD P_ISO W=1.435e-06 L=0.18e-06
M11 VDD A1 net_001 VDD P_ISO W=1.435e-06 L=0.18e-06
M12 net_001 A0 Q VDD P_ISO W=1.435e-06 L=0.18e-06
M13 net_001 A0 Q VDD P_ISO W=1.435e-06 L=0.18e-06
M14 Q A0 net_001 VDD P_ISO W=1.435e-06 L=0.18e-06
M15 VDD B0 Q VDD P_ISO W=1.435e-06 L=0.18e-06
M16 VDD B0 Q VDD P_ISO W=1.435e-06 L=0.18e-06
M17 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI21_X0_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_000 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_000 B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M3 VDD A1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M4 Q A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI21_X1_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 net_000 A1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_000 B0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VDD A1 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M4 Q A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI21_X2_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M4 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI21_X3_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M3 VSS A1 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M4 Q B0 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M5 Q B0 net_000 VSS N_ISO W=0.79e-06 L=0.18e-06
M6 VDD A1 net_001 VDD P_ISO W=0.865e-06 L=0.18e-06
M7 Q A0 net_001 VDD P_ISO W=0.865e-06 L=0.18e-06
M8 Q A0 net_002 VDD P_ISO W=0.865e-06 L=0.18e-06
M9 VDD A1 net_002 VDD P_ISO W=0.865e-06 L=0.18e-06
M10 VDD B0 Q VDD P_ISO W=0.865e-06 L=0.18e-06
M11 VDD B0 Q VDD P_ISO W=0.865e-06 L=0.18e-06
.ends

.subckt OAI21_X4_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI21_X6_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_000 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI21_X8_18_SVT_WB A0 A1 B0 Q VDD VSS
*.PININFO A0:I A1:I B0:I Q:O VDD:B VSS:B
M0 VSS A1 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M1 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A0 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M6 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_000 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI221_X0_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 net_000 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_001 C0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q A1 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_001 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q B0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD C0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M8 VDD A1 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q A0 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI221_X1_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 net_000 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 C0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q A1 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_001 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q B0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD C0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD A1 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q A0 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI221_X2_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 C0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD B1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI221_X4_18_SVT_WB A0 A1 B0 B1 C0 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I Q:O VDD:B VSS:B
M0 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_001 C0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_001 C0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_001 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD C0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD A1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q A0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI222_X0_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 VSS C1 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS C0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 B0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_001 B1 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 Q A1 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_001 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VDD C1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q C0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_003 B0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 VDD A1 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 Q A0 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI222_X1_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 VSS C1 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS C0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_001 B0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_001 B1 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q A1 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_001 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VDD C1 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q C0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_003 B0 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 VDD A1 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 Q A0 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI222_X2_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 VSS C1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_000 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD C1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q C0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_004 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI222_X4_18_SVT_WB A0 A1 B0 B1 C0 C1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I C0:I C1:I Q:O VDD:B VSS:B
M0 VSS C0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS C0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 B0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_001 B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_000 B1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_001 B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_001 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q A1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 Q A0 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 Q C0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD C1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD C1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q C0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD B1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD B1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q B0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q A0 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD A1 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD A1 net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 Q A0 net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI22_X0_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 B0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_000 A1 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD B1 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q B0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q A0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD A1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI22_X1_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_000 B0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q A0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_000 A1 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VDD B1 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 Q B0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 Q A0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD A1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI22_X2_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD B1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 Q B0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_002 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI22_X4_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD B1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q B0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B1 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q A0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI22_X8_18_SVT_WB A0 A1 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_001 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 net_002 VSS N_ISO W=0.715e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_001 B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_004 A0 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A1 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_001 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 net_002 VDD P_ISO W=0.815e-06 L=0.18e-06
M16 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI31_X0_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 net_000 A2 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_000 A0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_000 B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VDD A2 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_002 A1 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 Q A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI31_X1_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 net_000 A2 VSS VSS N_ISO W=0.575e-06 L=0.18e-06
M1 net_000 A1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_000 A0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_000 B0 Q VSS N_ISO W=0.575e-06 L=0.18e-06
M4 VDD A2 net_001 VDD P_ISO W=0.525e-06 L=0.18e-06
M5 net_002 A1 net_001 VDD P_ISO W=0.525e-06 L=0.18e-06
M6 Q A0 net_002 VDD P_ISO W=0.525e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=0.525e-06 L=0.18e-06
.ends

.subckt OAI31_X2_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 VSS A2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_000 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VDD A2 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M5 net_002 A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_002 A0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI31_X4_18_SVT_WB A0 A1 A2 B0 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I Q:O VDD:B VSS:B
M0 VSS A2 net_000 VSS N_ISO W=0.71e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_000 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD A2 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_002 A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_004 A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD A2 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B0 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI32_X0_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 A2 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 A1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_000 B0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_000 B1 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD A2 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 net_002 A1 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q A0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI32_X1_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 net_000 A2 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_000 A1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_000 B0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_000 B1 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD A2 net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_002 A1 net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q A0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI32_X2_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VDD A2 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_002 A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q B0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI32_X4_18_SVT_WB A0 A1 A2 B0 B1 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I Q:O VDD:B VSS:B
M0 VSS A2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS A2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 B0 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD A2 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_002 A1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q A0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_004 A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD A2 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q B0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q B0 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD B1 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI33_X0_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 net_000 B2 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 net_000 B1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_000 B0 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_000 A0 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_000 A1 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_000 A2 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VDD B2 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_002 B1 net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q B0 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M10 net_004 A1 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD A2 net_004 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt OAI33_X1_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 net_000 B2 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 net_000 B1 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_000 B0 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_000 A0 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_000 A1 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_000 A2 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VDD B2 net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_002 B1 net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 Q B0 net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 net_004 A1 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 VDD A2 net_004 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OAI33_X2_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 VSS B2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 A1 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A2 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VDD B2 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_002 B1 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q B0 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q A0 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_004 A1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A2 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OAI33_X4_18_SVT_WB A0 A1 A2 B0 B1 B2 Q VDD VSS
*.PININFO A0:I A1:I A2:I B0:I B1:I B2:I Q:O VDD:B VSS:B
M0 VSS B2 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B1 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A0 net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_000 A1 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A2 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD B2 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_004 B1 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_001 B0 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_001 A0 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_006 A1 net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD A2 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR2_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_0 A Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M4 VDD B net_0 VDD P_ISO W=0.42e-06 L=0.18e-06
M5 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OR2_X12_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q_neg B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_0_2 A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B net_0_2 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_0_1 B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 Q_neg A net_0_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_0_0 A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD B net_0_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M20 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_0 A Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M4 VDD B net_0 VDD P_ISO W=0.575e-06 L=0.18e-06
M5 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0 A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M5 VDD B net_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR2_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q_neg B VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M1 VSS A Q_neg VSS N_ISO W=0.785e-06 L=0.18e-06
M2 Q_neg A VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M3 VSS B Q_neg VSS N_ISO W=0.785e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_0_1 B VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M8 Q_neg A net_0_1 VDD P_ISO W=0.86e-06 L=0.18e-06
M9 net_0_0 A Q_neg VDD P_ISO W=0.86e-06 L=0.18e-06
M10 VDD B net_0_0 VDD P_ISO W=0.86e-06 L=0.18e-06
M11 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 Q_neg B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_0_1 B VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q_neg A net_0_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_0_0 A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_0_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M14 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR3_X1_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M1 Q_neg B VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS C Q_neg VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_0 A Q_neg VDD P_ISO W=0.42e-06 L=0.18e-06
M5 net_1 B net_0 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD C net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OR3_X12_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 Q net_000 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M15 net_002 A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_000 A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_003 A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_004 B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD C net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD C net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_002 B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_006 B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD C net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M28 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M29 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR3_X2_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M1 Q_neg B VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS C Q_neg VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_0 A Q_neg VDD P_ISO W=0.575e-06 L=0.18e-06
M5 net_1 B net_0 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD C net_1 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR3_X4_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M1 Q_neg B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_0 A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_1 B net_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD C net_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR3_X6_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 Q_neg C VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M1 VSS B Q_neg VSS N_ISO W=0.785e-06 L=0.18e-06
M2 Q_neg A VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M3 VSS A Q_neg VSS N_ISO W=0.785e-06 L=0.18e-06
M4 Q_neg B VSS VSS N_ISO W=0.785e-06 L=0.18e-06
M5 VSS C Q_neg VSS N_ISO W=0.785e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_1_1 C VDD VDD P_ISO W=0.86e-06 L=0.18e-06
M10 net_0_1 B net_1_1 VDD P_ISO W=0.86e-06 L=0.18e-06
M11 Q_neg A net_0_1 VDD P_ISO W=0.86e-06 L=0.18e-06
M12 net_0_0 A Q_neg VDD P_ISO W=0.86e-06 L=0.18e-06
M13 net_1_0 B net_0_0 VDD P_ISO W=0.86e-06 L=0.18e-06
M14 VDD C net_1_0 VDD P_ISO W=0.86e-06 L=0.18e-06
M15 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR3_X8_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 Q_neg C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M2 Q_neg A VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M4 Q_neg B VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS C Q_neg VSS N_ISO W=1.05e-06 L=0.18e-06
M6 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q Q_neg VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS Q_neg Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_1_1 C VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_0_1 B net_1_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 Q_neg A net_0_1 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_0_0 A Q_neg VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_1_0 B net_0_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD C net_1_0 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q Q_neg VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD Q_neg Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR4_X1_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.425e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.425e-06 L=0.18e-06
M2 VSS C net_000 VSS N_ISO W=0.425e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=0.425e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_000 A net_001 VDD P_ISO W=0.475e-06 L=0.18e-06
M6 net_002 B net_001 VDD P_ISO W=0.475e-06 L=0.18e-06
M7 net_003 C net_002 VDD P_ISO W=0.475e-06 L=0.18e-06
M8 VDD D net_003 VDD P_ISO W=0.475e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt OR4_X12_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_000 C VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD D net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_002 C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_003 B net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_003 A net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_000 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_005 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 net_005 C net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD D net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR4_X2_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS C net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 net_002 B net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_003 C net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_003 D VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR4_X4_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 net_000 A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 net_002 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_003 C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR4_X6_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_000 A net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_002 B net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 net_003 C net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD D net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt OR4_X8_18_SVT_WB A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:B VSS:B
M0 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS A net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS C net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS D net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD D net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_002 C net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_002 B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_000 A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_000 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_004 B net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_006 C net_005 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD D net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_000 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFQN_X1_18_SVT_WB D SE SI CK QN VDD VSS
*.PININFO D:I SE:I SI:I CK:I QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.83e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_009 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 VSS net_009 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M16 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M17 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M19 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M23 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M24 net_006 net_000 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_008 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_006 net_008 VDD P_ISO W=0.59e-06 L=0.18e-06
M27 net_009 net_000 net_008 VDD P_ISO W=0.67e-06 L=0.18e-06
M28 net_009 net_005 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M29 VDD net_011 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 VDD net_009 net_011 VDD P_ISO W=0.415e-06 L=0.18e-06
M31 VDD net_009 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFQN_X2_18_SVT_WB D SE SI CK QN VDD VSS
*.PININFO D:I SE:I SI:I CK:I QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.83e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_009 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 VSS net_009 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M16 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M17 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M19 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M23 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M24 net_006 net_000 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_008 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_006 net_008 VDD P_ISO W=0.59e-06 L=0.18e-06
M27 net_009 net_000 net_008 VDD P_ISO W=0.67e-06 L=0.18e-06
M28 net_009 net_005 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M29 VDD net_011 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 VDD net_009 net_011 VDD P_ISO W=0.415e-06 L=0.18e-06
M31 VDD net_009 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFQN_X4_18_SVT_WB D SE SI CK QN VDD VSS
*.PININFO D:I SE:I SI:I CK:I QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.83e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_009 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 VSS net_009 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M16 VSS net_009 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M18 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M24 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M25 net_006 net_000 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_008 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_006 net_008 VDD P_ISO W=0.59e-06 L=0.18e-06
M28 net_009 net_000 net_008 VDD P_ISO W=0.67e-06 L=0.18e-06
M29 net_009 net_005 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 VDD net_011 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M31 VDD net_009 net_011 VDD P_ISO W=0.415e-06 L=0.18e-06
M32 VDD net_009 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_009 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFQ_X1_18_SVT_WB D SE SI CK Q VDD VSS
*.PININFO D:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.83e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_009 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 VSS net_011 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M16 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M17 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M19 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M23 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M24 net_006 net_000 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_008 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_006 net_008 VDD P_ISO W=0.72e-06 L=0.18e-06
M27 net_008 net_000 net_009 VDD P_ISO W=0.67e-06 L=0.18e-06
M28 net_009 net_005 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M29 VDD net_011 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 VDD net_009 net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M31 VDD net_011 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFQ_X2_18_SVT_WB D SE SI CK Q VDD VSS
*.PININFO D:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.83e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 net_000 net_009 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 net_011 VSS N_ISO W=0.625e-06 L=0.18e-06
M15 VSS net_011 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M16 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M17 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M19 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M23 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M24 net_006 net_000 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M25 VDD net_008 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_006 net_008 VDD P_ISO W=0.72e-06 L=0.18e-06
M27 net_008 net_000 net_009 VDD P_ISO W=0.67e-06 L=0.18e-06
M28 net_009 net_005 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M29 VDD net_011 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 VDD net_009 net_011 VDD P_ISO W=0.59e-06 L=0.18e-06
M31 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFQ_X4_18_SVT_WB D SE SI CK Q VDD VSS
*.PININFO D:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.83e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_009 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 net_011 VSS N_ISO W=0.625e-06 L=0.18e-06
M15 VSS net_011 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M16 VSS net_011 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M18 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M24 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M25 net_006 net_000 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD net_008 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_006 net_008 VDD P_ISO W=0.72e-06 L=0.18e-06
M28 net_008 net_000 net_009 VDD P_ISO W=0.67e-06 L=0.18e-06
M29 net_009 net_005 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 VDD net_011 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M31 VDD net_009 net_011 VDD P_ISO W=0.59e-06 L=0.18e-06
M32 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFQ_X8_18_SVT_WB D SE SI CK Q VDD VSS
*.PININFO D:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.245e-06 L=0.18e-06
M10 net_008 net_006 VSS VSS N_ISO W=0.83e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 net_000 net_009 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 net_011 VSS N_ISO W=0.625e-06 L=0.18e-06
M15 VSS net_011 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M16 VSS net_011 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M17 VSS net_011 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M18 VSS net_011 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M27 net_006 net_000 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_008 net_014 VDD P_ISO W=0.22e-06 L=0.18e-06
M29 VDD net_006 net_008 VDD P_ISO W=0.72e-06 L=0.18e-06
M30 net_008 net_000 net_009 VDD P_ISO W=0.67e-06 L=0.18e-06
M31 net_009 net_005 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M32 VDD net_011 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M33 VDD net_009 net_011 VDD P_ISO W=0.59e-06 L=0.18e-06
M34 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFRQ_X1_18_SVT_WB D RN SE SI CK Q VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 net_008 RN net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.825e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_010 net_000 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_013 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M15 VSS RN net_012 VSS N_ISO W=0.42e-06 L=0.18e-06
M16 net_013 net_010 net_012 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M18 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M19 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M25 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M26 net_016 net_000 net_006 VDD P_ISO W=0.425e-06 L=0.18e-06
M27 VDD RN net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M28 VDD net_009 net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M29 VDD net_006 net_009 VDD P_ISO W=0.72e-06 L=0.18e-06
M30 net_010 net_000 net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M31 net_010 net_005 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M32 VDD net_013 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M33 VDD RN net_013 VDD P_ISO W=0.415e-06 L=0.18e-06
M34 VDD net_010 net_013 VDD P_ISO W=0.455e-06 L=0.18e-06
M35 VDD net_013 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFRQ_X2_18_SVT_WB D RN SE SI CK Q VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 net_008 RN net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.825e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_010 net_000 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_013 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M15 VSS RN net_012 VSS N_ISO W=0.53e-06 L=0.18e-06
M16 net_013 net_010 net_012 VSS N_ISO W=0.53e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M18 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M19 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M25 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M26 net_016 net_000 net_006 VDD P_ISO W=0.425e-06 L=0.18e-06
M27 VDD RN net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M28 VDD net_009 net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M29 VDD net_006 net_009 VDD P_ISO W=0.72e-06 L=0.18e-06
M30 net_010 net_000 net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M31 net_010 net_005 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M32 VDD net_013 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M33 VDD RN net_013 VDD P_ISO W=0.415e-06 L=0.18e-06
M34 VDD net_010 net_013 VDD P_ISO W=0.715e-06 L=0.18e-06
M35 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFRQ_X4_18_SVT_WB D RN SE SI CK Q VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 net_008 RN net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.825e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_010 net_000 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_013 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M15 VSS RN net_012 VSS N_ISO W=0.53e-06 L=0.18e-06
M16 net_013 net_010 net_012 VSS N_ISO W=0.53e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M18 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M27 net_016 net_000 net_006 VDD P_ISO W=0.425e-06 L=0.18e-06
M28 VDD RN net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M29 VDD net_009 net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M30 VDD net_006 net_009 VDD P_ISO W=0.72e-06 L=0.18e-06
M31 net_010 net_000 net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M32 net_010 net_005 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M33 VDD net_013 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M34 VDD RN net_013 VDD P_ISO W=0.415e-06 L=0.18e-06
M35 VDD net_010 net_013 VDD P_ISO W=0.715e-06 L=0.18e-06
M36 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFRQ_X8_18_SVT_WB D RN SE SI CK Q VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 net_008 RN net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 net_009 net_006 VSS VSS N_ISO W=0.825e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_010 net_000 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_013 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M15 VSS RN net_012 VSS N_ISO W=0.53e-06 L=0.18e-06
M16 net_013 net_010 net_012 VSS N_ISO W=0.53e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M18 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M19 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M20 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M21 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M22 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M24 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M25 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M28 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M29 net_016 net_000 net_006 VDD P_ISO W=0.425e-06 L=0.18e-06
M30 VDD RN net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M31 VDD net_009 net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M32 VDD net_006 net_009 VDD P_ISO W=0.72e-06 L=0.18e-06
M33 net_010 net_000 net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M34 net_010 net_005 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M35 VDD net_013 net_017 VDD P_ISO W=0.22e-06 L=0.18e-06
M36 VDD RN net_013 VDD P_ISO W=0.415e-06 L=0.18e-06
M37 VDD net_010 net_013 VDD P_ISO W=0.715e-06 L=0.18e-06
M38 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFR_X1_18_SVT_WB D RN SE SI CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.425e-06 L=0.18e-06
M9 net_008 RN net_007 VSS N_ISO W=0.425e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.425e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.825e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_013 net_011 VSS N_ISO W=0.82e-06 L=0.18e-06
M15 VSS RN net_012 VSS N_ISO W=0.42e-06 L=0.18e-06
M16 net_013 net_010 net_012 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M18 VSS net_011 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M27 net_016 net_000 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD RN net_016 VDD P_ISO W=0.685e-06 L=0.18e-06
M29 VDD net_009 net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M30 VDD net_006 net_009 VDD P_ISO W=0.94e-06 L=0.18e-06
M31 net_009 net_000 net_010 VDD P_ISO W=0.67e-06 L=0.18e-06
M32 net_011 net_005 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M33 VDD net_013 net_011 VDD P_ISO W=0.85e-06 L=0.18e-06
M34 VDD RN net_013 VDD P_ISO W=0.415e-06 L=0.18e-06
M35 VDD net_010 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M36 VDD net_013 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M37 VDD net_011 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFR_X2_18_SVT_WB D RN SE SI CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.425e-06 L=0.18e-06
M9 net_008 RN net_007 VSS N_ISO W=0.425e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.425e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.825e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_013 net_011 VSS N_ISO W=0.82e-06 L=0.18e-06
M15 VSS RN net_012 VSS N_ISO W=0.82e-06 L=0.18e-06
M16 net_013 net_010 net_012 VSS N_ISO W=0.82e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M18 VSS net_011 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M27 net_016 net_000 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD RN net_016 VDD P_ISO W=0.685e-06 L=0.18e-06
M29 VDD net_009 net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M30 VDD net_006 net_009 VDD P_ISO W=0.94e-06 L=0.18e-06
M31 net_009 net_000 net_010 VDD P_ISO W=0.67e-06 L=0.18e-06
M32 net_011 net_005 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M33 VDD net_013 net_011 VDD P_ISO W=0.85e-06 L=0.18e-06
M34 VDD RN net_013 VDD P_ISO W=0.415e-06 L=0.18e-06
M35 VDD net_010 net_013 VDD P_ISO W=0.715e-06 L=0.18e-06
M36 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_011 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFR_X4_18_SVT_WB D RN SE SI CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.425e-06 L=0.18e-06
M9 net_008 RN net_007 VSS N_ISO W=0.425e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.425e-06 L=0.18e-06
M11 net_009 net_006 VSS VSS N_ISO W=0.825e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_013 net_011 VSS N_ISO W=0.82e-06 L=0.18e-06
M15 VSS RN net_012 VSS N_ISO W=0.82e-06 L=0.18e-06
M16 net_013 net_010 net_012 VSS N_ISO W=0.82e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M18 VSS net_013 Q VSS N_ISO W=0.98e-06 L=0.18e-06
M19 VSS net_011 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M20 VSS net_011 QN VSS N_ISO W=0.98e-06 L=0.18e-06
M21 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M22 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M24 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M25 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M28 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M29 net_016 net_000 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD RN net_016 VDD P_ISO W=0.685e-06 L=0.18e-06
M31 VDD net_009 net_016 VDD P_ISO W=0.425e-06 L=0.18e-06
M32 VDD net_006 net_009 VDD P_ISO W=0.94e-06 L=0.18e-06
M33 net_009 net_000 net_010 VDD P_ISO W=0.67e-06 L=0.18e-06
M34 net_011 net_005 net_010 VDD P_ISO W=0.42e-06 L=0.18e-06
M35 VDD net_013 net_011 VDD P_ISO W=0.85e-06 L=0.18e-06
M36 VDD RN net_013 VDD P_ISO W=0.415e-06 L=0.18e-06
M37 VDD net_010 net_013 VDD P_ISO W=0.715e-06 L=0.18e-06
M38 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_011 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_011 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFSQ_X1_18_SVT_WB D SE SI SN CK Q VDD VSS
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_009 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M11 net_009 SN net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.565e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 net_011 SN net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M15 VSS net_013 net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M16 VSS net_010 net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M18 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M19 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_003 D net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_000 net_005 VDD P_ISO W=0.6e-06 L=0.18e-06
M25 net_006 net_005 net_003 VDD P_ISO W=0.57e-06 L=0.18e-06
M26 net_006 net_000 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_009 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_006 net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M29 VDD SN net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M30 net_010 net_000 net_009 VDD P_ISO W=0.565e-06 L=0.18e-06
M31 net_010 net_005 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M32 VDD SN net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M33 VDD net_013 net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M34 VDD net_010 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M35 VDD net_013 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFSQ_X2_18_SVT_WB D SE SI SN CK Q VDD VSS
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_009 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M11 net_009 SN net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.565e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 net_011 SN net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M15 VSS net_013 net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M16 VSS net_010 net_013 VSS N_ISO W=0.66e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M19 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_000 net_005 VDD P_ISO W=0.6e-06 L=0.18e-06
M25 net_006 net_005 net_003 VDD P_ISO W=0.57e-06 L=0.18e-06
M26 net_006 net_000 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M27 VDD net_009 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_006 net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M29 VDD SN net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M30 net_010 net_000 net_009 VDD P_ISO W=0.565e-06 L=0.18e-06
M31 net_010 net_005 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M32 VDD SN net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M33 VDD net_013 net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M34 VDD net_010 net_013 VDD P_ISO W=0.66e-06 L=0.18e-06
M35 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFSQ_X4_18_SVT_WB D SE SI SN CK Q VDD VSS
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_009 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M11 net_009 SN net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.565e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 net_011 SN net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M15 VSS net_013 net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M16 VSS net_010 net_013 VSS N_ISO W=0.995e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_014 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.57e-06 L=0.18e-06
M27 net_006 net_000 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_009 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M29 VDD net_006 net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M30 VDD SN net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M31 net_010 net_000 net_009 VDD P_ISO W=0.565e-06 L=0.18e-06
M32 net_010 net_005 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M33 VDD SN net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M34 VDD net_013 net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M35 VDD net_010 net_013 VDD P_ISO W=0.995e-06 L=0.18e-06
M36 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFSQ_X8_18_SVT_WB D SE SI SN CK Q VDD VSS
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_009 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M11 net_009 SN net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.565e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 net_011 SN net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M15 VSS net_013 net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M16 VSS net_010 net_013 VSS N_ISO W=0.995e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M22 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD SE net_014 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M25 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M28 net_006 net_005 net_003 VDD P_ISO W=0.57e-06 L=0.18e-06
M29 net_006 net_000 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD net_009 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M31 VDD net_006 net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M32 VDD SN net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M33 net_010 net_000 net_009 VDD P_ISO W=0.565e-06 L=0.18e-06
M34 net_010 net_005 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M35 VDD SN net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M36 VDD net_013 net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M37 VDD net_010 net_013 VDD P_ISO W=0.995e-06 L=0.18e-06
M38 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFSR_X1_18_SVT_WB D RN SE SI SN CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.7e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.335e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.335e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_003 net_000 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_008 net_010 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 VSS RN net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 SN net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_011 net_005 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M14 net_012 net_000 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 net_012 SN net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M16 VSS net_015 net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS RN net_014 VSS N_ISO W=0.42e-06 L=0.18e-06
M18 net_015 net_011 net_014 VSS N_ISO W=0.42e-06 L=0.18e-06
M19 VSS net_015 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M20 VSS net_012 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M21 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M22 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD SE net_016 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_016 D net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 net_017 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_001 net_017 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M28 net_006 net_005 net_003 VDD P_ISO W=0.555e-06 L=0.18e-06
M29 net_006 net_000 net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M30 VDD net_010 net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M31 VDD RN net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M32 VDD net_006 net_010 VDD P_ISO W=0.45e-06 L=0.18e-06
M33 VDD SN net_010 VDD P_ISO W=0.45e-06 L=0.18e-06
M34 net_010 net_000 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M35 net_011 net_005 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M36 VDD SN net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M37 VDD net_015 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M38 VDD RN net_015 VDD P_ISO W=0.45e-06 L=0.18e-06
M39 VDD net_011 net_015 VDD P_ISO W=0.45e-06 L=0.18e-06
M40 VDD net_015 Q VDD P_ISO W=0.7e-06 L=0.18e-06
M41 VDD net_012 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFSR_X2_18_SVT_WB D RN SE SI SN CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.7e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.335e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.335e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_003 net_000 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_008 net_010 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 VSS RN net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 SN net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_011 net_005 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M14 net_012 net_000 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 net_012 SN net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M16 VSS net_015 net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS RN net_014 VSS N_ISO W=0.42e-06 L=0.18e-06
M18 net_015 net_011 net_014 VSS N_ISO W=0.42e-06 L=0.18e-06
M19 Q net_015 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_012 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M22 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD SE net_016 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_016 D net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 net_017 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_001 net_017 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M28 net_006 net_005 net_003 VDD P_ISO W=0.585e-06 L=0.18e-06
M29 net_006 net_000 net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M30 VDD net_010 net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M31 VDD RN net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M32 VDD net_006 net_010 VDD P_ISO W=0.45e-06 L=0.18e-06
M33 VDD SN net_010 VDD P_ISO W=0.45e-06 L=0.18e-06
M34 net_010 net_000 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M35 net_011 net_005 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M36 VDD SN net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M37 VDD net_015 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M38 VDD RN net_015 VDD P_ISO W=0.45e-06 L=0.18e-06
M39 VDD net_011 net_015 VDD P_ISO W=0.45e-06 L=0.18e-06
M40 VDD net_015 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_012 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFSR_X4_18_SVT_WB D RN SE SI SN CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.7e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.335e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.335e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_003 net_000 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_008 net_010 net_007 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 VSS RN net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M11 VSS net_006 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 SN net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_011 net_005 net_010 VSS N_ISO W=0.42e-06 L=0.18e-06
M14 net_012 net_000 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M15 net_012 SN net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M16 VSS net_015 net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS RN net_014 VSS N_ISO W=0.42e-06 L=0.18e-06
M18 net_015 net_011 net_014 VSS N_ISO W=0.42e-06 L=0.18e-06
M19 VSS net_015 Q VSS N_ISO W=0.82e-06 L=0.18e-06
M20 VSS net_015 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS net_012 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VSS net_012 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M23 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M24 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD SE net_016 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 net_016 D net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 net_017 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M28 VDD net_001 net_017 VDD P_ISO W=0.42e-06 L=0.18e-06
M29 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M30 net_006 net_005 net_003 VDD P_ISO W=0.585e-06 L=0.18e-06
M31 net_006 net_000 net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M32 VDD net_010 net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M33 VDD RN net_018 VDD P_ISO W=0.45e-06 L=0.18e-06
M34 VDD net_006 net_010 VDD P_ISO W=0.45e-06 L=0.18e-06
M35 VDD SN net_010 VDD P_ISO W=0.45e-06 L=0.18e-06
M36 net_011 net_000 net_010 VDD P_ISO W=0.45e-06 L=0.18e-06
M37 net_011 net_005 net_012 VDD P_ISO W=0.45e-06 L=0.18e-06
M38 VDD SN net_012 VDD P_ISO W=0.625e-06 L=0.18e-06
M39 VDD net_015 net_012 VDD P_ISO W=0.625e-06 L=0.18e-06
M40 VDD RN net_015 VDD P_ISO W=0.45e-06 L=0.18e-06
M41 VDD net_011 net_015 VDD P_ISO W=0.45e-06 L=0.18e-06
M42 VDD net_015 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M43 VDD net_015 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M44 VDD net_012 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M45 VDD net_012 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFS_X1_18_SVT_WB D SE SI SN CK Q QN VDD VSS
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_009 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M11 net_009 SN net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.565e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 net_011 SN net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M15 VSS net_013 net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M16 VSS net_010 net_013 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M18 VSS net_011 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.6e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.57e-06 L=0.18e-06
M27 net_006 net_000 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_009 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M29 VDD net_006 net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M30 VDD SN net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M31 net_010 net_000 net_009 VDD P_ISO W=0.565e-06 L=0.18e-06
M32 net_010 net_005 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M33 VDD SN net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M34 VDD net_013 net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M35 VDD net_010 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M36 VDD net_013 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M37 VDD net_011 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFS_X2_18_SVT_WB D SE SI SN CK Q QN VDD VSS
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_009 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M11 net_009 SN net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.565e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 net_011 SN net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M15 VSS net_013 net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M16 VSS net_010 net_013 VSS N_ISO W=0.995e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_011 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_014 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.57e-06 L=0.18e-06
M27 net_006 net_000 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_009 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M29 VDD net_006 net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M30 VDD SN net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M31 net_010 net_000 net_009 VDD P_ISO W=0.565e-06 L=0.18e-06
M32 net_010 net_005 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M33 VDD SN net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M34 VDD net_013 net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M35 VDD net_010 net_013 VDD P_ISO W=0.995e-06 L=0.18e-06
M36 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_011 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFS_X4_18_SVT_WB D SE SI SN CK Q QN VDD VSS
*.PININFO D:I SE:I SI:I SN:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.585e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_009 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M11 net_009 SN net_008 VSS N_ISO W=0.935e-06 L=0.18e-06
M12 net_010 net_005 net_009 VSS N_ISO W=0.565e-06 L=0.18e-06
M13 net_011 net_000 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 net_011 SN net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M15 VSS net_013 net_012 VSS N_ISO W=0.655e-06 L=0.18e-06
M16 VSS net_010 net_013 VSS N_ISO W=0.995e-06 L=0.18e-06
M17 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_013 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_011 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_011 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M22 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD SE net_014 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 net_014 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M25 net_015 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M26 VDD net_001 net_015 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M28 net_006 net_005 net_003 VDD P_ISO W=0.57e-06 L=0.18e-06
M29 net_006 net_000 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD net_009 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M31 VDD net_006 net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M32 VDD SN net_009 VDD P_ISO W=0.64e-06 L=0.18e-06
M33 net_010 net_000 net_009 VDD P_ISO W=0.565e-06 L=0.18e-06
M34 net_010 net_005 net_011 VDD P_ISO W=0.45e-06 L=0.18e-06
M35 VDD SN net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M36 VDD net_013 net_011 VDD P_ISO W=0.655e-06 L=0.18e-06
M37 VDD net_010 net_013 VDD P_ISO W=0.995e-06 L=0.18e-06
M38 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_013 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M40 VDD net_011 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M41 VDD net_011 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFTR_X1_18_SVT_WB D RN SE SI CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS SI net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_004 RN net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS D net_004 VSS N_ISO W=0.815e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.61e-06 L=0.18e-06
M7 VSS net_005 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_007 net_005 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M9 net_007 net_006 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_007 net_009 VSS N_ISO W=0.585e-06 L=0.18e-06
M12 net_010 net_006 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_010 net_005 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_012 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M15 VSS net_010 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M16 VSS net_010 net_012 VSS N_ISO W=0.42e-06 L=0.18e-06
M17 VSS net_012 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M18 VDD SE net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD SI net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 net_002 net_000 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 net_014 SE net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD RN net_014 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD D net_014 VDD P_ISO W=0.915e-06 L=0.18e-06
M24 VDD CK net_005 VDD P_ISO W=0.435e-06 L=0.18e-06
M25 VDD net_005 net_006 VDD P_ISO W=0.725e-06 L=0.18e-06
M26 net_007 net_006 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 net_007 net_005 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_009 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M29 VDD net_007 net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 net_010 net_005 net_009 VDD P_ISO W=0.615e-06 L=0.18e-06
M31 net_010 net_006 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M32 VDD net_012 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M33 VDD net_010 QN VDD P_ISO W=0.575e-06 L=0.18e-06
M34 VDD net_010 net_012 VDD P_ISO W=0.42e-06 L=0.18e-06
M35 VDD net_012 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFFTR_X2_18_SVT_WB D RN SE SI CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS SI net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_004 RN net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS D net_004 VSS N_ISO W=0.815e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.61e-06 L=0.18e-06
M7 VSS net_005 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_007 net_005 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M9 net_007 net_006 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_007 net_009 VSS N_ISO W=0.585e-06 L=0.18e-06
M12 net_010 net_006 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_010 net_005 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_012 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M15 VSS net_010 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_010 net_012 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_012 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VDD SE net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD SI net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 net_002 net_000 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 net_014 SE net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD RN net_014 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD D net_014 VDD P_ISO W=0.915e-06 L=0.18e-06
M24 VDD CK net_005 VDD P_ISO W=0.435e-06 L=0.18e-06
M25 VDD net_005 net_006 VDD P_ISO W=0.725e-06 L=0.18e-06
M26 net_007 net_006 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M27 net_007 net_005 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD net_009 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M29 VDD net_007 net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M30 net_010 net_005 net_009 VDD P_ISO W=0.63e-06 L=0.18e-06
M31 net_010 net_006 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M32 VDD net_012 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M33 VDD net_010 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M34 VDD net_010 net_012 VDD P_ISO W=1.15e-06 L=0.18e-06
M35 VDD net_012 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFFTR_X4_18_SVT_WB D RN SE SI CK Q QN VDD VSS
*.PININFO D:I RN:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS SI net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_004 RN net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS D net_004 VSS N_ISO W=0.815e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.61e-06 L=0.18e-06
M7 VSS net_005 net_006 VSS N_ISO W=0.42e-06 L=0.18e-06
M8 net_007 net_005 net_002 VSS N_ISO W=0.425e-06 L=0.18e-06
M9 net_007 net_006 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_009 net_008 VSS N_ISO W=0.22e-06 L=0.18e-06
M11 VSS net_007 net_009 VSS N_ISO W=0.575e-06 L=0.18e-06
M12 net_010 net_006 net_009 VSS N_ISO W=0.42e-06 L=0.18e-06
M13 net_010 net_005 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_012 net_011 VSS N_ISO W=0.22e-06 L=0.18e-06
M15 VSS net_010 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_010 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_010 net_012 VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_012 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_012 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VDD SE net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SI net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 net_002 net_000 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 net_014 SE net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD RN net_014 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD D net_014 VDD P_ISO W=0.915e-06 L=0.18e-06
M26 VDD CK net_005 VDD P_ISO W=0.435e-06 L=0.18e-06
M27 VDD net_005 net_006 VDD P_ISO W=0.725e-06 L=0.18e-06
M28 net_007 net_006 net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M29 net_007 net_005 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD net_009 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M31 VDD net_007 net_009 VDD P_ISO W=0.42e-06 L=0.18e-06
M32 net_010 net_005 net_009 VDD P_ISO W=0.605e-06 L=0.18e-06
M33 net_010 net_006 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M34 VDD net_012 net_016 VDD P_ISO W=0.22e-06 L=0.18e-06
M35 VDD net_010 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_010 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_010 net_012 VDD P_ISO W=1.15e-06 L=0.18e-06
M38 VDD net_012 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M39 VDD net_012 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFF_X1_18_SVT_WB D SE SI CK Q QN VDD VSS
*.PININFO D:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.61e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 net_000 net_009 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M15 VSS net_009 net_011 VSS N_ISO W=0.42e-06 L=0.18e-06
M16 VSS net_011 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M18 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M24 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M25 net_006 net_000 net_014 VDD P_ISO W=0.445e-06 L=0.18e-06
M26 VDD net_008 net_014 VDD P_ISO W=0.445e-06 L=0.18e-06
M27 net_008 net_006 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M28 net_009 net_000 net_008 VDD P_ISO W=0.625e-06 L=0.18e-06
M29 net_009 net_005 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD net_011 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M31 VDD net_009 QN VDD P_ISO W=0.575e-06 L=0.18e-06
M32 VDD net_009 net_011 VDD P_ISO W=0.42e-06 L=0.18e-06
M33 VDD net_011 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt SDFF_X2_18_SVT_WB D SE SI CK Q QN VDD VSS
*.PININFO D:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.615e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 net_000 net_009 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_009 net_011 VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_011 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M18 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M20 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M21 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M22 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M23 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M24 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M25 net_006 net_000 net_014 VDD P_ISO W=0.445e-06 L=0.18e-06
M26 VDD net_008 net_014 VDD P_ISO W=0.445e-06 L=0.18e-06
M27 net_008 net_006 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M28 net_009 net_000 net_008 VDD P_ISO W=0.59e-06 L=0.18e-06
M29 net_009 net_005 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD net_011 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M31 VDD net_009 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M32 VDD net_009 net_011 VDD P_ISO W=1.15e-06 L=0.18e-06
M33 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt SDFF_X4_18_SVT_WB D SE SI CK Q QN VDD VSS
*.PININFO D:I SE:I SI:I CK:I Q:O QN:O VDD:B VSS:B
M0 VSS CK net_000 VSS N_ISO W=0.585e-06 L=0.18e-06
M1 VSS SE net_002 VSS N_ISO W=0.22e-06 L=0.18e-06
M2 VSS SE net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 SI net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 net_003 D net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M5 VSS net_001 net_004 VSS N_ISO W=0.825e-06 L=0.18e-06
M6 VSS net_000 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 net_006 net_000 net_003 VSS N_ISO W=0.425e-06 L=0.18e-06
M8 net_006 net_005 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M9 VSS net_008 net_007 VSS N_ISO W=0.22e-06 L=0.18e-06
M10 VSS net_006 net_008 VSS N_ISO W=0.62e-06 L=0.18e-06
M11 net_009 net_005 net_008 VSS N_ISO W=0.42e-06 L=0.18e-06
M12 net_010 net_000 net_009 VSS N_ISO W=0.22e-06 L=0.18e-06
M13 VSS net_011 net_010 VSS N_ISO W=0.22e-06 L=0.18e-06
M14 VSS net_009 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_009 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_009 net_011 VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_011 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_011 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VDD CK net_000 VDD P_ISO W=0.565e-06 L=0.18e-06
M20 VDD SE net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M21 VDD SE net_012 VDD P_ISO W=0.535e-06 L=0.18e-06
M22 net_012 D net_003 VDD P_ISO W=0.535e-06 L=0.18e-06
M23 net_013 SI net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M24 VDD net_001 net_013 VDD P_ISO W=0.42e-06 L=0.18e-06
M25 VDD net_000 net_005 VDD P_ISO W=0.555e-06 L=0.18e-06
M26 net_006 net_005 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M27 net_006 net_000 net_014 VDD P_ISO W=0.445e-06 L=0.18e-06
M28 VDD net_008 net_014 VDD P_ISO W=0.445e-06 L=0.18e-06
M29 net_008 net_006 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M30 net_009 net_000 net_008 VDD P_ISO W=0.605e-06 L=0.18e-06
M31 net_009 net_005 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M32 VDD net_011 net_015 VDD P_ISO W=0.22e-06 L=0.18e-06
M33 VDD net_009 QN VDD P_ISO W=1.125e-06 L=0.18e-06
M34 VDD net_009 QN VDD P_ISO W=1.125e-06 L=0.18e-06
M35 VDD net_009 net_011 VDD P_ISO W=1.15e-06 L=0.18e-06
M36 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M37 VDD net_011 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TIEH_18_SVT_WB Q VDD VSS
*.PININFO Q:O VDD:B VSS:B
M0 VSS net_000 net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VDD net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt TIEL_18_SVT_WB Q VDD VSS
*.PININFO Q:O VDD:B VSS:B
M0 VSS net_001 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VDD net_001 net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt TLATNCA_X12_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.605e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_006 CK net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 net_007 net_003 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 net_008 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M21 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M22 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M23 VDD net_001 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M24 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M26 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M27 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M28 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M29 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M30 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M31 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M32 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M33 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M34 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M35 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M36 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M37 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNCA_X16_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.605e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_006 CK net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_007 net_003 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M22 net_008 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M23 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M24 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 VDD net_001 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M26 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M27 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M29 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M30 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M31 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M32 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M33 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M34 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M35 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M36 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M37 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M38 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M39 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M40 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M41 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNCA_X2_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_006 CK net_007 VSS N_ISO W=0.38e-06 L=0.18e-06
M8 VSS net_003 net_007 VSS N_ISO W=0.44e-06 L=0.18e-06
M9 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M11 net_001 net_004 net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M12 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD CK net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 VDD CK net_006 VDD P_ISO W=0.375e-06 L=0.18e-06
M18 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNCA_X20_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.605e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_006 CK net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M23 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M24 net_008 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M26 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M27 VDD net_001 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M28 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M29 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M31 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M32 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M33 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M34 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M35 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M36 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M37 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M38 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M39 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M40 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M41 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M42 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M43 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M44 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M45 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNCA_X3_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_006 CK net_007 VSS N_ISO W=0.38e-06 L=0.18e-06
M8 VSS net_003 net_007 VSS N_ISO W=0.44e-06 L=0.18e-06
M9 VSS net_006 ECK VSS N_ISO W=0.79e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=0.79e-06 L=0.18e-06
M11 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M12 net_001 net_004 net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD CK net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 VDD CK net_006 VDD P_ISO W=0.375e-06 L=0.18e-06
M19 VDD net_003 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M20 VDD net_006 ECK VDD P_ISO W=0.875e-06 L=0.18e-06
M21 VDD net_006 ECK VDD P_ISO W=0.875e-06 L=0.18e-06
.ends

.subckt TLATNCA_X4_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_007 CK net_006 VSS N_ISO W=0.38e-06 L=0.18e-06
M8 VSS net_003 net_007 VSS N_ISO W=0.855e-06 L=0.18e-06
M9 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M12 net_008 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M18 VDD CK net_006 VDD P_ISO W=0.375e-06 L=0.18e-06
M19 VDD net_003 net_006 VDD P_ISO W=0.88e-06 L=0.18e-06
M20 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M21 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNCA_X6_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 net_008 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M19 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M20 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M21 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M22 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M23 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNCA_X8_18_SVT_WB CK E ECK VDD VSS
*.PININFO CK:I E:I ECK:O VDD:B VSS:B
M0 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M6 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M7 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 net_008 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_001 net_005 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD net_003 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 net_006 CK VDD VDD P_ISO W=1.145e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M22 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M23 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M24 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M25 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNSR_X1_18_SVT_WB D GN RN SN Q QN VDD VSS
*.PININFO D:I GN:I RN:I SN:I Q:O QN:O VDD:B VSS:B
M0 VSS GN net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS RN net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M2 net_002 D net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M3 net_003 net_000 net_002 VSS N_ISO W=0.295e-06 L=0.18e-06
M4 net_003 GN net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M5 net_005 net_007 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.295e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M9 VSS net_007 net_008 VSS N_ISO W=0.44e-06 L=0.18e-06
M10 VSS net_007 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M12 VDD GN net_000 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 VDD RN net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 VDD D net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_003 GN net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 net_003 net_000 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_007 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_003 net_007 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD SN net_007 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 VDD net_007 net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M21 VDD net_007 QN VDD P_ISO W=0.575e-06 L=0.18e-06
M22 VDD net_008 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt TLATNSR_X2_18_SVT_WB D GN RN SN Q QN VDD VSS
*.PININFO D:I GN:I RN:I SN:I Q:O QN:O VDD:B VSS:B
M0 VSS GN net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS RN net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M2 net_002 D net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M3 net_003 net_000 net_002 VSS N_ISO W=0.295e-06 L=0.18e-06
M4 net_003 GN net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M5 net_005 net_007 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.295e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.6e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.6e-06 L=0.18e-06
M9 VSS net_007 net_008 VSS N_ISO W=0.7e-06 L=0.18e-06
M10 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD GN net_000 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 VDD RN net_003 VDD P_ISO W=0.585e-06 L=0.18e-06
M14 VDD D net_009 VDD P_ISO W=0.585e-06 L=0.18e-06
M15 net_003 GN net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 net_003 net_000 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_007 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_003 net_007 VDD P_ISO W=0.53e-06 L=0.18e-06
M19 VDD SN net_007 VDD P_ISO W=0.53e-06 L=0.18e-06
M20 VDD net_007 net_008 VDD P_ISO W=0.8e-06 L=0.18e-06
M21 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TLATNSR_X4_18_SVT_WB D GN RN SN Q QN VDD VSS
*.PININFO D:I GN:I RN:I SN:I Q:O QN:O VDD:B VSS:B
M0 VSS GN net_000 VSS N_ISO W=0.745e-06 L=0.18e-06
M1 VSS RN net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M2 net_002 D net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M3 net_003 net_000 net_002 VSS N_ISO W=0.295e-06 L=0.18e-06
M4 net_003 GN net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M5 net_005 net_007 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.295e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.595e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.595e-06 L=0.18e-06
M9 VSS net_007 net_008 VSS N_ISO W=1e-06 L=0.18e-06
M10 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_008 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 Q net_008 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD GN net_000 VDD P_ISO W=0.875e-06 L=0.18e-06
M15 VDD RN net_003 VDD P_ISO W=0.61e-06 L=0.18e-06
M16 VDD D net_009 VDD P_ISO W=0.61e-06 L=0.18e-06
M17 net_003 GN net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 net_003 net_000 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD net_007 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 VDD net_003 net_007 VDD P_ISO W=0.525e-06 L=0.18e-06
M21 VDD SN net_007 VDD P_ISO W=0.525e-06 L=0.18e-06
M22 VDD net_007 net_008 VDD P_ISO W=1.09e-06 L=0.18e-06
M23 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q net_008 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X12_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.605e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_006 CK net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VDD SE net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M21 net_009 E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M22 net_009 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M23 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M24 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 VDD net_001 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M26 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M27 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M28 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M29 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M30 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M31 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M32 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M33 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M34 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M35 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M36 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M37 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M38 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M39 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X16_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.605e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_006 CK net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VDD SE net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M23 net_009 E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M24 net_009 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M26 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M27 VDD net_001 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M28 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M29 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M30 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M31 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M32 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M33 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M34 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M35 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M36 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M37 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M38 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M39 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M40 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M41 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M42 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M43 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X2_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.56e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=0.38e-06 L=0.18e-06
M9 VSS net_003 net_007 VSS N_ISO W=0.44e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD SE net_008 VDD P_ISO W=0.57e-06 L=0.18e-06
M12 net_009 E net_008 VDD P_ISO W=0.57e-06 L=0.18e-06
M13 net_009 net_004 net_001 VDD P_ISO W=0.57e-06 L=0.18e-06
M14 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M19 VDD CK net_006 VDD P_ISO W=0.375e-06 L=0.18e-06
M20 VDD net_003 net_006 VDD P_ISO W=0.44e-06 L=0.18e-06
M21 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X20_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.605e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_006 CK net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M15 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M16 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M17 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M18 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M19 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M20 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M21 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M22 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M23 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M24 VDD SE net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M25 net_009 E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M26 net_009 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M27 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M28 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M29 VDD net_001 net_003 VDD P_ISO W=0.685e-06 L=0.18e-06
M30 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M31 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M32 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M33 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M34 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M35 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M36 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M37 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M38 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M39 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M40 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M41 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M42 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M43 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M44 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M45 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M46 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M47 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X3_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=0.38e-06 L=0.18e-06
M9 VSS net_003 net_007 VSS N_ISO W=0.485e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=0.79e-06 L=0.18e-06
M11 VSS net_006 ECK VSS N_ISO W=0.79e-06 L=0.18e-06
M12 VDD SE net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 net_009 E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 net_009 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 net_006 CK VDD VDD P_ISO W=0.375e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=0.49e-06 L=0.18e-06
M22 VDD net_006 ECK VDD P_ISO W=0.865e-06 L=0.18e-06
M23 VDD net_006 ECK VDD P_ISO W=0.865e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X4_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=0.38e-06 L=0.18e-06
M9 VSS net_003 net_007 VSS N_ISO W=0.855e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD SE net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 net_009 E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 net_009 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M20 net_006 CK VDD VDD P_ISO W=0.375e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=0.88e-06 L=0.18e-06
M22 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M23 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X6_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD SE net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 net_009 E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_009 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M21 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M22 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M23 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M24 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M25 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATNTSCA_X8_18_SVT_WB CK E SE ECK VDD VSS
*.PININFO CK:I E:I SE:I ECK:O VDD:B VSS:B
M0 VSS SE net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS E net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_001 net_005 net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_001 net_004 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M4 VSS net_003 net_002 VSS N_ISO W=0.44e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_005 net_004 VSS N_ISO W=0.47e-06 L=0.18e-06
M7 VSS CK net_005 VSS N_ISO W=0.25e-06 L=0.18e-06
M8 net_007 CK net_006 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_003 net_007 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_006 ECK VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD SE net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_009 E net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 net_009 net_004 net_001 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 net_001 net_005 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_003 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD net_001 net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 VDD net_005 net_004 VDD P_ISO W=0.44e-06 L=0.18e-06
M21 VDD CK net_005 VDD P_ISO W=0.22e-06 L=0.18e-06
M22 VDD CK net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M23 VDD net_003 net_006 VDD P_ISO W=1.145e-06 L=0.18e-06
M24 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M25 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M26 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
M27 VDD net_006 ECK VDD P_ISO W=1.145e-06 L=0.18e-06
.ends

.subckt TLATN_X1_18_SVT_WB D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
M0 VSS GN net_000 VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_002 GN net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 VSS net_004 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_004 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M8 VDD GN net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M9 VDD D net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M10 net_002 GN net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M11 net_002 net_000 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M12 net_006 net_004 VDD VDD P_ISO W=0.22e-06 L=0.18e-06
M13 VDD net_002 net_004 VDD P_ISO W=0.625e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M15 VDD net_004 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt TLATN_X2_18_SVT_WB D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
M0 VSS GN net_000 VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_002 GN net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 VSS net_004 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD GN net_000 VDD P_ISO W=0.65e-06 L=0.18e-06
M9 VDD D net_005 VDD P_ISO W=0.435e-06 L=0.18e-06
M10 net_002 GN net_005 VDD P_ISO W=0.435e-06 L=0.18e-06
M11 net_002 net_000 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M12 VDD net_004 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M13 VDD net_002 net_004 VDD P_ISO W=0.625e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_004 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TLATN_X4_18_SVT_WB D GN Q QN VDD VSS
*.PININFO D:I GN:I Q:O QN:O VDD:B VSS:B
M0 VSS GN net_000 VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 net_000 net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_002 GN net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 VSS net_004 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.995e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_004 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M9 QN net_004 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD GN net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M11 VDD D net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M12 net_002 GN net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 net_002 net_000 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M14 VDD net_004 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M15 VDD net_002 net_004 VDD P_ISO W=1.02e-06 L=0.18e-06
M16 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_004 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M19 QN net_004 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TLATSR_X1_18_SVT_WB D G RN SN Q QN VDD VSS
*.PININFO D:I G:I RN:I SN:I Q:O QN:O VDD:B VSS:B
M0 VSS G net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS RN net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M2 net_002 D net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M3 net_003 G net_002 VSS N_ISO W=0.295e-06 L=0.18e-06
M4 net_003 net_000 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M5 net_005 net_007 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.295e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M9 VSS net_007 net_008 VSS N_ISO W=0.44e-06 L=0.18e-06
M10 VSS net_007 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M12 VDD G net_000 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 VDD RN net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 VDD D net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_003 net_000 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 net_003 G net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_007 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_003 net_007 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD SN net_007 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 VDD net_007 net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M21 VDD net_007 QN VDD P_ISO W=0.575e-06 L=0.18e-06
M22 VDD net_008 Q VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt TLATSR_X2_18_SVT_WB D G RN SN Q QN VDD VSS
*.PININFO D:I G:I RN:I SN:I Q:O QN:O VDD:B VSS:B
M0 VSS G net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS RN net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M2 net_002 D net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M3 net_003 G net_002 VSS N_ISO W=0.295e-06 L=0.18e-06
M4 net_003 net_000 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M5 net_005 net_007 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.295e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M9 VSS net_007 net_008 VSS N_ISO W=0.44e-06 L=0.18e-06
M10 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_008 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VDD G net_000 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 VDD RN net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M14 VDD D net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 net_003 net_000 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 net_003 G net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 VDD net_007 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 VDD net_003 net_007 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD SN net_007 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 VDD net_007 net_008 VDD P_ISO W=0.44e-06 L=0.18e-06
M21 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TLATSR_X4_18_SVT_WB D G RN SN Q QN VDD VSS
*.PININFO D:I G:I RN:I SN:I Q:O QN:O VDD:B VSS:B
M0 VSS G net_000 VSS N_ISO W=0.44e-06 L=0.18e-06
M1 VSS RN net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M2 net_002 D net_001 VSS N_ISO W=0.295e-06 L=0.18e-06
M3 net_003 G net_002 VSS N_ISO W=0.295e-06 L=0.18e-06
M4 net_003 net_000 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M5 net_005 net_007 net_004 VSS N_ISO W=0.295e-06 L=0.18e-06
M6 VSS RN net_005 VSS N_ISO W=0.295e-06 L=0.18e-06
M7 VSS net_003 net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M8 net_007 SN net_006 VSS N_ISO W=0.5e-06 L=0.18e-06
M9 VSS net_007 net_008 VSS N_ISO W=1e-06 L=0.18e-06
M10 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_007 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_008 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 Q net_008 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M14 VDD G net_000 VDD P_ISO W=0.44e-06 L=0.18e-06
M15 VDD RN net_003 VDD P_ISO W=0.44e-06 L=0.18e-06
M16 VDD D net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M17 net_003 net_000 net_009 VDD P_ISO W=0.44e-06 L=0.18e-06
M18 net_003 G net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M19 VDD net_007 net_010 VDD P_ISO W=0.44e-06 L=0.18e-06
M20 net_007 net_003 VDD VDD P_ISO W=0.44e-06 L=0.18e-06
M21 VDD SN net_007 VDD P_ISO W=0.44e-06 L=0.18e-06
M22 VDD net_007 net_008 VDD P_ISO W=1.09e-06 L=0.18e-06
M23 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_007 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_008 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 Q net_008 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TLAT_X1_18_SVT_WB D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
M0 VSS G net_000 VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 G net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 VSS net_004 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_004 QN VSS N_ISO W=0.525e-06 L=0.18e-06
M8 VDD G net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M9 VDD D net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M10 net_002 net_000 net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M11 net_002 G net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M12 net_006 net_004 VDD VDD P_ISO W=0.22e-06 L=0.18e-06
M13 VDD net_002 net_004 VDD P_ISO W=0.625e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M15 VDD net_004 QN VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt TLAT_X2_18_SVT_WB D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
M0 VSS G net_000 VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 G net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 VSS net_004 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.44e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_004 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VDD G net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M9 VDD D net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M10 net_002 net_000 net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M11 net_002 G net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M12 VDD net_004 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M13 VDD net_002 net_004 VDD P_ISO W=0.625e-06 L=0.18e-06
M14 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_004 QN VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt TLAT_X4_18_SVT_WB D G Q QN VDD VSS
*.PININFO D:I G:I Q:O QN:O VDD:B VSS:B
M0 VSS G net_000 VSS N_ISO W=0.5e-06 L=0.18e-06
M1 VSS D net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M2 net_002 G net_001 VSS N_ISO W=0.44e-06 L=0.18e-06
M3 net_002 net_000 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M4 VSS net_004 net_003 VSS N_ISO W=0.22e-06 L=0.18e-06
M5 VSS net_002 net_004 VSS N_ISO W=0.995e-06 L=0.18e-06
M6 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_002 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_004 QN VSS N_ISO W=1.05e-06 L=0.18e-06
M9 QN net_004 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VDD G net_000 VDD P_ISO W=0.655e-06 L=0.18e-06
M11 VDD D net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M12 net_002 net_000 net_005 VDD P_ISO W=0.44e-06 L=0.18e-06
M13 net_002 G net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M14 VDD net_004 net_006 VDD P_ISO W=0.22e-06 L=0.18e-06
M15 VDD net_002 net_004 VDD P_ISO W=1.02e-06 L=0.18e-06
M16 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_002 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 VDD net_004 QN VDD P_ISO W=1.15e-06 L=0.18e-06
M19 QN net_004 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR2PG_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q A net_001 VSS N_ISO W=0.9e-06 L=0.18e-06
M4 net_000 net_002 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M5 VDD B net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD net_000 net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD A net_002 VDD P_ISO W=0.725e-06 L=0.18e-06
M8 net_000 A Q VDD P_ISO W=1.3e-06 L=0.18e-06
M9 net_001 net_002 Q VDD P_ISO W=1.3e-06 L=0.18e-06
.ends

.subckt XNOR2PG_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS net_000 net_001 VSS N_ISO W=0.9e-06 L=0.18e-06
M2 VSS A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q A net_001 VSS N_ISO W=0.9e-06 L=0.18e-06
M4 net_000 net_002 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M5 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M7 VDD A net_002 VDD P_ISO W=0.725e-06 L=0.18e-06
M8 net_000 A Q VDD P_ISO W=1.3e-06 L=0.18e-06
M9 net_001 net_002 Q VDD P_ISO W=1.3e-06 L=0.18e-06
.ends

.subckt XNOR2PG_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 net_001 net_000 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS net_000 net_001 VSS N_ISO W=0.9e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 Q A net_001 VSS N_ISO W=0.9e-06 L=0.18e-06
M6 net_000 net_002 Q VSS N_ISO W=0.9e-06 L=0.18e-06
M7 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD A net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M12 net_000 A Q VDD P_ISO W=1.3e-06 L=0.18e-06
M13 Q net_002 net_001 VDD P_ISO W=1.3e-06 L=0.18e-06
.ends

.subckt XNOR2PG_X6_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B net_000 VSS N_ISO W=0.88e-06 L=0.18e-06
M3 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M4 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M5 Q A net_001 VSS N_ISO W=0.88e-06 L=0.18e-06
M6 net_001 A Q VSS N_ISO W=0.88e-06 L=0.18e-06
M7 VSS A net_002 VSS N_ISO W=0.88e-06 L=0.18e-06
M8 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M15 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M16 Q A net_000 VDD P_ISO W=1.32e-06 L=0.18e-06
M17 net_000 A Q VDD P_ISO W=1.32e-06 L=0.18e-06
M18 VDD A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR2PG_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M2 VSS B net_000 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 VSS B net_000 VSS N_ISO W=0.88e-06 L=0.18e-06
M4 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M5 net_000 net_002 Q VSS N_ISO W=0.88e-06 L=0.18e-06
M6 Q A net_001 VSS N_ISO W=0.88e-06 L=0.18e-06
M7 net_001 A Q VSS N_ISO W=0.88e-06 L=0.18e-06
M8 VSS A net_002 VSS N_ISO W=0.88e-06 L=0.18e-06
M9 VSS net_000 net_001 VSS N_ISO W=0.88e-06 L=0.18e-06
M10 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M18 net_001 net_002 Q VDD P_ISO W=1.32e-06 L=0.18e-06
M19 Q A net_000 VDD P_ISO W=1.32e-06 L=0.18e-06
M20 Q A net_000 VDD P_ISO W=1.32e-06 L=0.18e-06
M21 VDD A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_000 net_001 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR2_X0_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_001 A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 net_002 net_000 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 Q A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_002 B Q VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VDD A net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q net_000 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 net_003 A Q VDD P_ISO W=0.42e-06 L=0.18e-06
M9 VDD B net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt XNOR2_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 Q B net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD A net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 Q net_000 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_003 A Q VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD B net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt XNOR2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_2 A x1 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_2 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 net_1 x1 VSS VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A net_1 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_1 B Q VSS N_ISO W=1.05e-06 L=0.18e-06
M5 x1 A VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B x1 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 Q x1 VDD VDD P_ISO W=1.15e-06 L=0.18e-06
M8 net_0 A Q VDD P_ISO W=1.15e-06 L=0.18e-06
M9 VDD B net_0 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 net_003 A net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD B net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_001 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 net_001 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_003 A net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 VDD B net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 VDD net_000 net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_001 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 net_001 B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR3_X0_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_004 net_001 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS C net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 VSS net_003 net_005 VSS N_ISO W=0.755e-06 L=0.18e-06
M8 Q net_001 net_005 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 net_005 C Q VSS N_ISO W=0.42e-06 L=0.18e-06
M10 net_006 A net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD B net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD net_000 net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M13 net_007 A net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M14 net_007 B net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M15 net_003 net_001 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M16 VDD C net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M18 net_008 net_001 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M19 VDD C net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt XNOR3_X1_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 net_002 B VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_003 net_001 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS C net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 VSS net_003 net_005 VSS N_ISO W=0.525e-06 L=0.18e-06
M8 net_005 net_001 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M9 Q C net_005 VSS N_ISO W=0.525e-06 L=0.18e-06
M10 net_006 A net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD B net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD net_000 net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M13 net_001 A net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M14 net_007 B net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M15 net_003 net_001 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M16 VDD C net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M18 net_008 net_001 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M19 VDD C net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt XNOR3_X2_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 A net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 net_002 B VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_003 net_001 net_004 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VSS C net_004 VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_003 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 Q net_001 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 Q C net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_000 A net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD B net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD net_000 net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 net_001 A net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M14 net_001 B net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M15 net_003 net_001 VDD VDD P_ISO W=0.575e-06 L=0.18e-06
M16 VDD C net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_008 net_001 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD C net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR3_X4_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VSS C net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_003 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_004 net_001 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS C net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_000 A net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD B net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M14 VDD net_000 net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_001 A net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_001 B net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_008 net_001 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M18 VDD C net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M19 VDD net_003 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 net_004 net_001 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 net_004 C net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XNOR3_X8_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VSS C net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_003 net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_004 net_001 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS C net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_004 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_000 A net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M15 VDD B net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M16 VDD net_000 net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_001 A net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_001 B net_007 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 net_008 net_001 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M20 VDD C net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M21 VDD net_003 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_004 net_001 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 net_004 C net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_004 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XOR2NG_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS net_002 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q net_000 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 B Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VDD B net_000 VDD P_ISO W=0.555e-06 L=0.18e-06
M6 net_000 net_002 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M7 net_002 net_000 Q VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD A net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt XOR2NG_X1P5_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS net_002 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 Q net_000 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 Q B net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS A net_002 VSS N_ISO W=0.71e-06 L=0.18e-06
M5 VDD B net_000 VDD P_ISO W=1.15e-06 L=0.18e-06
M6 net_000 net_002 Q VDD P_ISO W=0.665e-06 L=0.18e-06
M7 net_002 net_000 Q VDD P_ISO W=0.665e-06 L=0.18e-06
M8 VDD A net_002 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XOR2_X0_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 x1 A VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B x1 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q x1 VSS VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_0 A Q VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS B net_0 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 net_2 A x1 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B net_2 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 net_1 x1 VDD VDD P_ISO W=0.42e-06 L=0.18e-06
M8 Q A net_1 VDD P_ISO W=0.42e-06 L=0.18e-06
M9 net_1 B Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt XOR2_X1_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 Q net_000 VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_001 A Q VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 net_000 A net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M6 VDD B net_002 VDD P_ISO W=0.42e-06 L=0.18e-06
M7 VDD net_000 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 net_003 A Q VDD P_ISO W=0.575e-06 L=0.18e-06
M9 Q B net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt XOR2_X2_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M3 Q A net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_000 A net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M6 VDD B net_002 VDD P_ISO W=0.575e-06 L=0.18e-06
M7 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M8 Q A net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M9 Q B net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XOR2_X3_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_003 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_003 Q VSS N_ISO W=0.785e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=0.785e-06 L=0.18e-06
M7 VDD A net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD B net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_003 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_003 Q VDD P_ISO W=0.86e-06 L=0.18e-06
M13 VDD net_003 Q VDD P_ISO W=0.86e-06 L=0.18e-06
.ends

.subckt XOR2_X4_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_003 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VDD A net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M8 VDD B net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M9 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M10 net_003 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M11 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XOR2_X8_18_SVT_WB A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:B VSS:B
M0 net_000 A net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_003 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 net_003 B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M6 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VDD A net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M10 VDD B net_000 VDD P_ISO W=0.575e-06 L=0.18e-06
M11 VDD net_000 net_003 VDD P_ISO W=1.15e-06 L=0.18e-06
M12 net_003 A net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M13 VDD B net_004 VDD P_ISO W=1.15e-06 L=0.18e-06
M14 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M15 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M16 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_003 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XOR3_X0_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_001 A net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS C net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=0.42e-06 L=0.18e-06
M8 Q net_001 net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M9 VSS C net_004 VSS N_ISO W=0.42e-06 L=0.18e-06
M10 net_005 A net_000 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD B net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD net_000 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M13 net_006 A net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M14 net_006 B net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M15 net_007 net_001 net_003 VDD P_ISO W=0.42e-06 L=0.18e-06
M16 VDD C net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 VDD net_003 net_008 VDD P_ISO W=0.42e-06 L=0.18e-06
M18 net_008 net_001 Q VDD P_ISO W=0.42e-06 L=0.18e-06
M19 net_008 C Q VDD P_ISO W=0.42e-06 L=0.18e-06
.ends

.subckt XOR3_X1_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M3 net_002 A net_001 VSS N_ISO W=0.42e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=0.42e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M6 VSS C net_003 VSS N_ISO W=0.42e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=0.525e-06 L=0.18e-06
M8 Q net_001 net_004 VSS N_ISO W=0.525e-06 L=0.18e-06
M9 VSS C net_004 VSS N_ISO W=0.525e-06 L=0.18e-06
M10 net_000 A net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD B net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD net_000 net_006 VDD P_ISO W=0.42e-06 L=0.18e-06
M13 net_006 A net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M14 net_006 B net_001 VDD P_ISO W=0.42e-06 L=0.18e-06
M15 net_003 net_001 net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M16 VDD C net_007 VDD P_ISO W=0.42e-06 L=0.18e-06
M17 VDD net_003 net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M18 Q net_001 net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
M19 Q C net_008 VDD P_ISO W=0.575e-06 L=0.18e-06
.ends

.subckt XOR3_X2_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.42e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M3 net_002 A net_001 VSS N_ISO W=0.525e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=0.525e-06 L=0.18e-06
M5 VSS net_001 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VSS C net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_003 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_004 net_001 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M9 VSS C net_004 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 net_000 A net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M11 VDD B net_005 VDD P_ISO W=0.42e-06 L=0.18e-06
M12 VDD net_000 net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 net_006 A net_001 VDD P_ISO W=0.575e-06 L=0.18e-06
M14 net_001 B net_006 VDD P_ISO W=0.575e-06 L=0.18e-06
M15 net_007 net_001 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M16 VDD C net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M17 VDD net_003 net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 Q net_001 net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 Q C net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XOR3_X4_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_003 net_001 net_004 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 VSS C net_004 VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_003 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_006 net_001 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_006 C net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_006 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_006 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 net_000 A net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M13 VDD B net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M14 VDD net_000 net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M15 net_001 A net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M16 net_001 B net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 VDD net_001 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M18 VDD C net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M19 VDD net_003 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M20 net_006 net_001 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M21 VDD C net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 VDD net_006 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD net_006 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.subckt XOR3_X8_18_SVT_WB A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:B VSS:B
M0 VSS A net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M1 VSS B net_000 VSS N_ISO W=0.525e-06 L=0.18e-06
M2 VSS net_000 net_001 VSS N_ISO W=1.05e-06 L=0.18e-06
M3 net_001 A net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M4 VSS B net_002 VSS N_ISO W=1.05e-06 L=0.18e-06
M5 net_004 net_001 net_003 VSS N_ISO W=0.525e-06 L=0.18e-06
M6 net_004 C VSS VSS N_ISO W=0.525e-06 L=0.18e-06
M7 VSS net_003 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M8 net_006 net_001 net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M9 net_006 C net_005 VSS N_ISO W=1.05e-06 L=0.18e-06
M10 VSS net_006 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M11 VSS net_006 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M12 VSS net_006 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M13 VSS net_006 Q VSS N_ISO W=1.05e-06 L=0.18e-06
M14 net_000 A net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M15 VDD B net_007 VDD P_ISO W=0.575e-06 L=0.18e-06
M16 VDD net_000 net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M17 net_001 A net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M18 net_001 B net_008 VDD P_ISO W=1.15e-06 L=0.18e-06
M19 VDD net_001 net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M20 VDD C net_003 VDD P_ISO W=0.575e-06 L=0.18e-06
M21 VDD net_003 net_006 VDD P_ISO W=1.15e-06 L=0.18e-06
M22 net_006 net_001 net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M23 VDD C net_009 VDD P_ISO W=1.15e-06 L=0.18e-06
M24 VDD net_006 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M25 VDD net_006 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M26 VDD net_006 Q VDD P_ISO W=1.15e-06 L=0.18e-06
M27 VDD net_006 Q VDD P_ISO W=1.15e-06 L=0.18e-06
.ends

.option scale = 1e-6
